
module betterNeighborsInMyCluster_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_inc_3 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module betterNeighborsInMyCluster_DW01_add_11 ( A, B, CI, SUM, CO );
  input [17:0] A;
  input [17:0] B;
  output [17:0] SUM;
  input CI;
  output CO;
  wire   \A[2] , \A[1] , \A[0] , n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66;
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX0 U2 ( .INP(n38), .ZN(n14) );
  INVX0 U3 ( .INP(n35), .ZN(n13) );
  INVX0 U4 ( .INP(n31), .ZN(n12) );
  INVX0 U5 ( .INP(n19), .ZN(n9) );
  INVX0 U6 ( .INP(n65), .ZN(n8) );
  INVX0 U7 ( .INP(n27), .ZN(n11) );
  INVX0 U8 ( .INP(n59), .ZN(n7) );
  INVX0 U9 ( .INP(n23), .ZN(n10) );
  INVX0 U10 ( .INP(n56), .ZN(n6) );
  AND2X1 U11 ( .IN1(A[3]), .IN2(B[3]), .Q(n1) );
  INVX0 U12 ( .INP(n43), .ZN(n3) );
  OAI21X1 U13 ( .IN1(n39), .IN2(n40), .IN3(n41), .QN(SUM[17]) );
  INVX0 U14 ( .INP(n39), .ZN(n15) );
  INVX0 U15 ( .INP(n52), .ZN(n5) );
  INVX0 U16 ( .INP(n47), .ZN(n4) );
  XOR2X1 U17 ( .IN1(A[3]), .IN2(B[3]), .Q(SUM[3]) );
  XNOR2X1 U18 ( .IN1(n16), .IN2(n17), .Q(SUM[9]) );
  NOR2X0 U19 ( .IN1(n9), .IN2(n18), .QN(n17) );
  XOR2X1 U20 ( .IN1(n20), .IN2(n21), .Q(SUM[8]) );
  NAND2X0 U21 ( .IN1(n10), .IN2(n22), .QN(n20) );
  XOR2X1 U22 ( .IN1(n24), .IN2(n25), .Q(SUM[7]) );
  NAND2X0 U23 ( .IN1(n11), .IN2(n26), .QN(n24) );
  XNOR2X1 U24 ( .IN1(n28), .IN2(n29), .Q(SUM[6]) );
  NOR2X0 U25 ( .IN1(n12), .IN2(n30), .QN(n29) );
  XNOR2X1 U26 ( .IN1(n32), .IN2(n33), .Q(SUM[5]) );
  NOR2X0 U27 ( .IN1(n13), .IN2(n34), .QN(n33) );
  XOR2X1 U28 ( .IN1(n1), .IN2(n36), .Q(SUM[4]) );
  NOR2X0 U29 ( .IN1(n37), .IN2(n38), .QN(n36) );
  XOR2X1 U30 ( .IN1(n42), .IN2(n40), .Q(SUM[16]) );
  OA21X1 U31 ( .IN1(n43), .IN2(n44), .IN3(n45), .Q(n40) );
  NAND2X0 U32 ( .IN1(n15), .IN2(n41), .QN(n42) );
  NAND2X0 U33 ( .IN1(B[16]), .IN2(A[16]), .QN(n41) );
  NOR2X0 U34 ( .IN1(B[16]), .IN2(A[16]), .QN(n39) );
  XOR2X1 U35 ( .IN1(n46), .IN2(n44), .Q(SUM[15]) );
  OA21X1 U36 ( .IN1(n47), .IN2(n48), .IN3(n49), .Q(n44) );
  NAND2X0 U37 ( .IN1(n3), .IN2(n45), .QN(n46) );
  NAND2X0 U38 ( .IN1(B[15]), .IN2(A[15]), .QN(n45) );
  NOR2X0 U39 ( .IN1(B[15]), .IN2(A[15]), .QN(n43) );
  XOR2X1 U40 ( .IN1(n50), .IN2(n48), .Q(SUM[14]) );
  OA21X1 U41 ( .IN1(n51), .IN2(n52), .IN3(n53), .Q(n48) );
  NAND2X0 U42 ( .IN1(n4), .IN2(n49), .QN(n50) );
  NAND2X0 U43 ( .IN1(B[14]), .IN2(A[14]), .QN(n49) );
  NOR2X0 U44 ( .IN1(B[14]), .IN2(A[14]), .QN(n47) );
  XOR2X1 U45 ( .IN1(n54), .IN2(n51), .Q(SUM[13]) );
  OA21X1 U46 ( .IN1(n55), .IN2(n56), .IN3(n57), .Q(n51) );
  NAND2X0 U47 ( .IN1(n5), .IN2(n53), .QN(n54) );
  NAND2X0 U48 ( .IN1(B[13]), .IN2(A[13]), .QN(n53) );
  NOR2X0 U49 ( .IN1(B[13]), .IN2(A[13]), .QN(n52) );
  XOR2X1 U50 ( .IN1(n58), .IN2(n55), .Q(SUM[12]) );
  OA21X1 U51 ( .IN1(n59), .IN2(n60), .IN3(n61), .Q(n55) );
  NAND2X0 U52 ( .IN1(n6), .IN2(n57), .QN(n58) );
  NAND2X0 U53 ( .IN1(B[12]), .IN2(A[12]), .QN(n57) );
  NOR2X0 U54 ( .IN1(B[12]), .IN2(A[12]), .QN(n56) );
  XOR2X1 U55 ( .IN1(n62), .IN2(n60), .Q(SUM[11]) );
  OA21X1 U56 ( .IN1(n63), .IN2(n64), .IN3(n65), .Q(n60) );
  NAND2X0 U57 ( .IN1(n7), .IN2(n61), .QN(n62) );
  NAND2X0 U58 ( .IN1(B[11]), .IN2(A[11]), .QN(n61) );
  NOR2X0 U59 ( .IN1(B[11]), .IN2(A[11]), .QN(n59) );
  XNOR2X1 U60 ( .IN1(n64), .IN2(n66), .Q(SUM[10]) );
  NOR2X0 U61 ( .IN1(n8), .IN2(n63), .QN(n66) );
  NOR2X0 U62 ( .IN1(B[10]), .IN2(A[10]), .QN(n63) );
  NAND2X0 U63 ( .IN1(B[10]), .IN2(A[10]), .QN(n65) );
  OA21X1 U64 ( .IN1(n18), .IN2(n16), .IN3(n19), .Q(n64) );
  NAND2X0 U65 ( .IN1(B[9]), .IN2(A[9]), .QN(n19) );
  OA21X1 U66 ( .IN1(n21), .IN2(n23), .IN3(n22), .Q(n16) );
  NAND2X0 U67 ( .IN1(B[8]), .IN2(A[8]), .QN(n22) );
  NOR2X0 U68 ( .IN1(B[8]), .IN2(A[8]), .QN(n23) );
  OA21X1 U69 ( .IN1(n27), .IN2(n25), .IN3(n26), .Q(n21) );
  NAND2X0 U70 ( .IN1(B[7]), .IN2(A[7]), .QN(n26) );
  OA21X1 U71 ( .IN1(n30), .IN2(n28), .IN3(n31), .Q(n25) );
  NAND2X0 U72 ( .IN1(B[6]), .IN2(A[6]), .QN(n31) );
  OA21X1 U73 ( .IN1(n32), .IN2(n34), .IN3(n35), .Q(n28) );
  NAND2X0 U74 ( .IN1(B[5]), .IN2(A[5]), .QN(n35) );
  NOR2X0 U75 ( .IN1(B[5]), .IN2(A[5]), .QN(n34) );
  AOI21X1 U76 ( .IN1(n14), .IN2(n1), .IN3(n37), .QN(n32) );
  AND2X1 U77 ( .IN1(B[4]), .IN2(A[4]), .Q(n37) );
  NOR2X0 U78 ( .IN1(B[4]), .IN2(A[4]), .QN(n38) );
  NOR2X0 U79 ( .IN1(B[6]), .IN2(A[6]), .QN(n30) );
  NOR2X0 U80 ( .IN1(B[7]), .IN2(A[7]), .QN(n27) );
  NOR2X0 U81 ( .IN1(B[9]), .IN2(A[9]), .QN(n18) );
endmodule


module betterNeighborsInMyCluster_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [3:0] A;
  input [15:0] B;
  output [19:0] PRODUCT;
  input TC;
  wire   \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] , \ab[3][11] ,
         \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] , \ab[3][6] ,
         \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] , \ab[3][1] ,
         \ab[3][0] , \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[3][0] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] ,
         \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] ,
         \A1[3] , \A1[2] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30;
  assign \ab[3][15]  = B[15];
  assign \ab[3][14]  = B[14];
  assign \ab[3][13]  = B[13];
  assign \ab[3][12]  = B[12];
  assign \ab[3][11]  = B[11];
  assign \ab[3][10]  = B[10];
  assign \ab[3][9]  = B[9];
  assign \ab[3][8]  = B[8];
  assign \ab[3][7]  = B[7];
  assign \ab[3][6]  = B[6];
  assign \ab[3][5]  = B[5];
  assign \ab[3][4]  = B[4];
  assign \ab[3][3]  = B[3];
  assign \ab[3][2]  = B[2];
  assign \ab[3][1]  = B[1];
  assign PRODUCT[1] = \ab[3][0] ;
  assign \ab[3][0]  = B[0];

  betterNeighborsInMyCluster_DW01_add_11 FS_1 ( .A({1'b0, \ab[3][15] , 
        \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , 
        \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \SUMB[3][0] , \ab[3][1] }), .B({1'b0, n30, n14, n15, n13, n12, n7, n6, 
        n5, n4, n10, n9, n8, n11, n3, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(
        PRODUCT[19:2]) );
  AND2X1 U2 ( .IN1(n21), .IN2(\SUMB[3][1] ), .Q(n3) );
  AND2X1 U3 ( .IN1(n19), .IN2(\SUMB[3][6] ), .Q(n4) );
  AND2X1 U4 ( .IN1(n20), .IN2(\SUMB[3][7] ), .Q(n5) );
  AND2X1 U5 ( .IN1(n24), .IN2(\SUMB[3][8] ), .Q(n6) );
  AND2X1 U6 ( .IN1(n25), .IN2(\SUMB[3][9] ), .Q(n7) );
  AND2X1 U7 ( .IN1(n16), .IN2(\SUMB[3][3] ), .Q(n8) );
  AND2X1 U8 ( .IN1(n17), .IN2(\SUMB[3][4] ), .Q(n9) );
  AND2X1 U9 ( .IN1(n18), .IN2(\SUMB[3][5] ), .Q(n10) );
  AND2X1 U10 ( .IN1(n22), .IN2(\SUMB[3][2] ), .Q(n11) );
  AND2X1 U11 ( .IN1(n23), .IN2(\SUMB[3][10] ), .Q(n12) );
  AND2X1 U12 ( .IN1(n27), .IN2(\SUMB[3][11] ), .Q(n13) );
  AND2X1 U13 ( .IN1(n29), .IN2(\SUMB[3][13] ), .Q(n14) );
  AND2X1 U14 ( .IN1(n28), .IN2(\SUMB[3][12] ), .Q(n15) );
  AND2X1 U15 ( .IN1(\ab[3][2] ), .IN2(\ab[3][4] ), .Q(n16) );
  AND2X1 U16 ( .IN1(\ab[3][3] ), .IN2(\ab[3][5] ), .Q(n17) );
  AND2X1 U17 ( .IN1(\ab[3][4] ), .IN2(\ab[3][6] ), .Q(n18) );
  AND2X1 U18 ( .IN1(\ab[3][5] ), .IN2(\ab[3][7] ), .Q(n19) );
  AND2X1 U19 ( .IN1(\ab[3][6] ), .IN2(\ab[3][8] ), .Q(n20) );
  AND2X1 U20 ( .IN1(\ab[3][0] ), .IN2(\ab[3][2] ), .Q(n21) );
  AND2X1 U21 ( .IN1(\ab[3][1] ), .IN2(\ab[3][3] ), .Q(n22) );
  AND2X1 U22 ( .IN1(\ab[3][9] ), .IN2(\ab[3][11] ), .Q(n23) );
  AND2X1 U23 ( .IN1(\ab[3][7] ), .IN2(\ab[3][9] ), .Q(n24) );
  AND2X1 U24 ( .IN1(\ab[3][8] ), .IN2(\ab[3][10] ), .Q(n25) );
  AND2X1 U25 ( .IN1(\ab[3][13] ), .IN2(\ab[3][15] ), .Q(n26) );
  AND2X1 U26 ( .IN1(\ab[3][10] ), .IN2(\ab[3][12] ), .Q(n27) );
  AND2X1 U27 ( .IN1(\ab[3][11] ), .IN2(\ab[3][13] ), .Q(n28) );
  AND2X1 U28 ( .IN1(\ab[3][12] ), .IN2(\ab[3][14] ), .Q(n29) );
  AND2X1 U29 ( .IN1(n26), .IN2(\ab[3][14] ), .Q(n30) );
  XOR2X1 U30 ( .IN1(n21), .IN2(\SUMB[3][1] ), .Q(\A1[2] ) );
  XOR2X1 U31 ( .IN1(n22), .IN2(\SUMB[3][2] ), .Q(\A1[3] ) );
  XOR2X1 U32 ( .IN1(n16), .IN2(\SUMB[3][3] ), .Q(\A1[4] ) );
  XOR2X1 U33 ( .IN1(n17), .IN2(\SUMB[3][4] ), .Q(\A1[5] ) );
  XOR2X1 U34 ( .IN1(n18), .IN2(\SUMB[3][5] ), .Q(\A1[6] ) );
  XOR2X1 U35 ( .IN1(n19), .IN2(\SUMB[3][6] ), .Q(\A1[7] ) );
  XOR2X1 U36 ( .IN1(n20), .IN2(\SUMB[3][7] ), .Q(\A1[8] ) );
  XOR2X1 U37 ( .IN1(n24), .IN2(\SUMB[3][8] ), .Q(\A1[9] ) );
  XOR2X1 U38 ( .IN1(n25), .IN2(\SUMB[3][9] ), .Q(\A1[10] ) );
  XOR2X1 U39 ( .IN1(n23), .IN2(\SUMB[3][10] ), .Q(\A1[11] ) );
  XOR2X1 U40 ( .IN1(n27), .IN2(\SUMB[3][11] ), .Q(\A1[12] ) );
  XOR2X1 U41 ( .IN1(n29), .IN2(\SUMB[3][13] ), .Q(\A1[14] ) );
  XOR2X1 U42 ( .IN1(n26), .IN2(\ab[3][14] ), .Q(\A1[15] ) );
  XOR2X1 U43 ( .IN1(n28), .IN2(\SUMB[3][12] ), .Q(\A1[13] ) );
  XOR2X1 U44 ( .IN1(\ab[3][2] ), .IN2(\ab[3][0] ), .Q(\SUMB[3][0] ) );
  XOR2X1 U45 ( .IN1(\ab[3][3] ), .IN2(\ab[3][1] ), .Q(\SUMB[3][1] ) );
  XOR2X1 U46 ( .IN1(\ab[3][4] ), .IN2(\ab[3][2] ), .Q(\SUMB[3][2] ) );
  XOR2X1 U47 ( .IN1(\ab[3][5] ), .IN2(\ab[3][3] ), .Q(\SUMB[3][3] ) );
  XOR2X1 U48 ( .IN1(\ab[3][6] ), .IN2(\ab[3][4] ), .Q(\SUMB[3][4] ) );
  XOR2X1 U49 ( .IN1(\ab[3][7] ), .IN2(\ab[3][5] ), .Q(\SUMB[3][5] ) );
  XOR2X1 U50 ( .IN1(\ab[3][8] ), .IN2(\ab[3][6] ), .Q(\SUMB[3][6] ) );
  XOR2X1 U51 ( .IN1(\ab[3][9] ), .IN2(\ab[3][7] ), .Q(\SUMB[3][7] ) );
  XOR2X1 U52 ( .IN1(\ab[3][10] ), .IN2(\ab[3][8] ), .Q(\SUMB[3][8] ) );
  XOR2X1 U53 ( .IN1(\ab[3][11] ), .IN2(\ab[3][9] ), .Q(\SUMB[3][9] ) );
  XOR2X1 U54 ( .IN1(\ab[3][12] ), .IN2(\ab[3][10] ), .Q(\SUMB[3][10] ) );
  XOR2X1 U55 ( .IN1(\ab[3][13] ), .IN2(\ab[3][11] ), .Q(\SUMB[3][11] ) );
  XOR2X1 U56 ( .IN1(\ab[3][14] ), .IN2(\ab[3][12] ), .Q(\SUMB[3][12] ) );
  XOR2X1 U57 ( .IN1(\ab[3][15] ), .IN2(\ab[3][13] ), .Q(\SUMB[3][13] ) );
endmodule


module betterNeighborsInMyCluster_DW01_add_10 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] ,
         \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n3,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62;
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  INVX0 U2 ( .INP(n56), .ZN(n12) );
  INVX0 U3 ( .INP(n52), .ZN(n11) );
  INVX0 U4 ( .INP(n44), .ZN(n9) );
  INVX0 U5 ( .INP(n48), .ZN(n10) );
  INVX0 U6 ( .INP(n40), .ZN(n8) );
  INVX0 U7 ( .INP(n32), .ZN(n6) );
  INVX0 U8 ( .INP(n36), .ZN(n7) );
  INVX0 U9 ( .INP(n28), .ZN(n5) );
  INVX0 U10 ( .INP(n24), .ZN(n4) );
  INVX0 U11 ( .INP(n20), .ZN(n3) );
  INVX0 U12 ( .INP(n60), .ZN(n13) );
  AND2X1 U13 ( .IN1(n59), .IN2(n1), .Q(SUM[15]) );
  OR2X1 U14 ( .IN1(B[15]), .IN2(A[15]), .Q(n1) );
  INVX0 U15 ( .INP(n15), .ZN(n2) );
  XNOR3X1 U16 ( .IN1(B[28]), .IN2(A[28]), .IN3(n14), .Q(SUM[28]) );
  OA21X1 U17 ( .IN1(n15), .IN2(n16), .IN3(n17), .Q(n14) );
  XOR2X1 U18 ( .IN1(n18), .IN2(n16), .Q(SUM[27]) );
  OA21X1 U19 ( .IN1(n19), .IN2(n20), .IN3(n21), .Q(n16) );
  NAND2X0 U20 ( .IN1(n2), .IN2(n17), .QN(n18) );
  NAND2X0 U21 ( .IN1(B[27]), .IN2(A[27]), .QN(n17) );
  NOR2X0 U22 ( .IN1(B[27]), .IN2(A[27]), .QN(n15) );
  XOR2X1 U23 ( .IN1(n22), .IN2(n19), .Q(SUM[26]) );
  OA21X1 U24 ( .IN1(n23), .IN2(n24), .IN3(n25), .Q(n19) );
  NAND2X0 U25 ( .IN1(n3), .IN2(n21), .QN(n22) );
  NAND2X0 U26 ( .IN1(B[26]), .IN2(A[26]), .QN(n21) );
  NOR2X0 U27 ( .IN1(B[26]), .IN2(A[26]), .QN(n20) );
  XOR2X1 U28 ( .IN1(n26), .IN2(n23), .Q(SUM[25]) );
  OA21X1 U29 ( .IN1(n27), .IN2(n28), .IN3(n29), .Q(n23) );
  NAND2X0 U30 ( .IN1(n4), .IN2(n25), .QN(n26) );
  NAND2X0 U31 ( .IN1(B[25]), .IN2(A[25]), .QN(n25) );
  NOR2X0 U32 ( .IN1(B[25]), .IN2(A[25]), .QN(n24) );
  XOR2X1 U33 ( .IN1(n30), .IN2(n27), .Q(SUM[24]) );
  OA21X1 U34 ( .IN1(n31), .IN2(n32), .IN3(n33), .Q(n27) );
  NAND2X0 U35 ( .IN1(n5), .IN2(n29), .QN(n30) );
  NAND2X0 U36 ( .IN1(B[24]), .IN2(A[24]), .QN(n29) );
  NOR2X0 U37 ( .IN1(B[24]), .IN2(A[24]), .QN(n28) );
  XOR2X1 U38 ( .IN1(n34), .IN2(n31), .Q(SUM[23]) );
  OA21X1 U39 ( .IN1(n35), .IN2(n36), .IN3(n37), .Q(n31) );
  NAND2X0 U40 ( .IN1(n6), .IN2(n33), .QN(n34) );
  NAND2X0 U41 ( .IN1(B[23]), .IN2(A[23]), .QN(n33) );
  NOR2X0 U42 ( .IN1(B[23]), .IN2(A[23]), .QN(n32) );
  XOR2X1 U43 ( .IN1(n38), .IN2(n35), .Q(SUM[22]) );
  OA21X1 U44 ( .IN1(n39), .IN2(n40), .IN3(n41), .Q(n35) );
  NAND2X0 U45 ( .IN1(n7), .IN2(n37), .QN(n38) );
  NAND2X0 U46 ( .IN1(B[22]), .IN2(A[22]), .QN(n37) );
  NOR2X0 U47 ( .IN1(B[22]), .IN2(A[22]), .QN(n36) );
  XOR2X1 U48 ( .IN1(n42), .IN2(n39), .Q(SUM[21]) );
  OA21X1 U49 ( .IN1(n43), .IN2(n44), .IN3(n45), .Q(n39) );
  NAND2X0 U50 ( .IN1(n8), .IN2(n41), .QN(n42) );
  NAND2X0 U51 ( .IN1(B[21]), .IN2(A[21]), .QN(n41) );
  NOR2X0 U52 ( .IN1(B[21]), .IN2(A[21]), .QN(n40) );
  XOR2X1 U53 ( .IN1(n46), .IN2(n43), .Q(SUM[20]) );
  OA21X1 U54 ( .IN1(n47), .IN2(n48), .IN3(n49), .Q(n43) );
  NAND2X0 U55 ( .IN1(n9), .IN2(n45), .QN(n46) );
  NAND2X0 U56 ( .IN1(B[20]), .IN2(A[20]), .QN(n45) );
  NOR2X0 U57 ( .IN1(B[20]), .IN2(A[20]), .QN(n44) );
  XOR2X1 U58 ( .IN1(n50), .IN2(n47), .Q(SUM[19]) );
  OA21X1 U59 ( .IN1(n51), .IN2(n52), .IN3(n53), .Q(n47) );
  NAND2X0 U60 ( .IN1(n10), .IN2(n49), .QN(n50) );
  NAND2X0 U61 ( .IN1(B[19]), .IN2(A[19]), .QN(n49) );
  NOR2X0 U62 ( .IN1(B[19]), .IN2(A[19]), .QN(n48) );
  XOR2X1 U63 ( .IN1(n54), .IN2(n51), .Q(SUM[18]) );
  OA21X1 U64 ( .IN1(n55), .IN2(n56), .IN3(n57), .Q(n51) );
  NAND2X0 U65 ( .IN1(n11), .IN2(n53), .QN(n54) );
  NAND2X0 U66 ( .IN1(B[18]), .IN2(A[18]), .QN(n53) );
  NOR2X0 U67 ( .IN1(B[18]), .IN2(A[18]), .QN(n52) );
  XOR2X1 U68 ( .IN1(n58), .IN2(n55), .Q(SUM[17]) );
  OA21X1 U69 ( .IN1(n59), .IN2(n60), .IN3(n61), .Q(n55) );
  NAND2X0 U70 ( .IN1(n12), .IN2(n57), .QN(n58) );
  NAND2X0 U71 ( .IN1(B[17]), .IN2(A[17]), .QN(n57) );
  NOR2X0 U72 ( .IN1(B[17]), .IN2(A[17]), .QN(n56) );
  XOR2X1 U73 ( .IN1(n62), .IN2(n59), .Q(SUM[16]) );
  NAND2X0 U74 ( .IN1(n13), .IN2(n61), .QN(n62) );
  NAND2X0 U75 ( .IN1(B[16]), .IN2(A[16]), .QN(n61) );
  NOR2X0 U76 ( .IN1(B[16]), .IN2(A[16]), .QN(n60) );
  NAND2X0 U77 ( .IN1(B[15]), .IN2(A[15]), .QN(n59) );
endmodule


module betterNeighborsInMyCluster_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][15] , \ab[15][14] , \ab[15][13] , \ab[15][12] , \ab[15][11] ,
         \ab[15][10] , \ab[15][9] , \ab[15][8] , \ab[15][7] , \ab[15][6] ,
         \ab[15][5] , \ab[15][4] , \ab[15][3] , \ab[15][2] , \ab[15][1] ,
         \ab[15][0] , \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] ,
         \ab[14][11] , \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] ,
         \ab[14][6] , \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] ,
         \ab[14][1] , \ab[14][0] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][15] ,
         \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] , \ab[11][10] ,
         \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] , \ab[11][5] ,
         \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] , \ab[11][0] ,
         \ab[10][15] , \ab[10][14] , \ab[10][13] , \ab[10][12] , \ab[10][11] ,
         \ab[10][10] , \ab[10][9] , \ab[10][8] , \ab[10][7] , \ab[10][6] ,
         \ab[10][5] , \ab[10][4] , \ab[10][3] , \ab[10][2] , \ab[10][1] ,
         \ab[10][0] , \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] ,
         \ab[9][11] , \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] ,
         \ab[9][6] , \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] ,
         \ab[9][1] , \ab[9][0] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][15] ,
         \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] , \ab[6][10] ,
         \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] , \ab[6][5] ,
         \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] , \ab[6][0] ,
         \ab[5][15] , \ab[5][14] , \ab[5][13] , \ab[5][12] , \ab[5][11] ,
         \ab[5][10] , \ab[5][9] , \ab[5][8] , \ab[5][7] , \ab[5][6] ,
         \ab[5][5] , \ab[5][4] , \ab[5][3] , \ab[5][2] , \ab[5][1] ,
         \ab[5][0] , \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] ,
         \ab[4][11] , \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] ,
         \ab[4][6] , \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] ,
         \ab[4][1] , \ab[4][0] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][15] , \ab[2][14] ,
         \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] ,
         \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] ,
         \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][15] ,
         \ab[1][14] , \ab[1][13] , \ab[1][12] , \ab[1][11] , \ab[1][10] ,
         \ab[1][9] , \ab[1][8] , \ab[1][7] , \ab[1][6] , \ab[1][5] ,
         \ab[1][4] , \ab[1][3] , \ab[1][2] , \ab[1][1] , \ab[1][0] ,
         \ab[0][15] , \ab[0][14] , \ab[0][13] , \ab[0][12] , \ab[0][11] ,
         \ab[0][10] , \ab[0][9] , \ab[0][8] , \ab[0][7] , \ab[0][6] ,
         \ab[0][5] , \ab[0][4] , \ab[0][3] , \ab[0][2] , \ab[0][1] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][14] , \CARRYB[14][13] , \CARRYB[14][12] ,
         \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] , \CARRYB[14][8] ,
         \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[14][0] ,
         \CARRYB[13][14] , \CARRYB[13][13] , \CARRYB[13][12] ,
         \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] ,
         \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] , \CARRYB[13][4] ,
         \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] , \CARRYB[13][0] ,
         \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] , \CARRYB[12][4] ,
         \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[12][0] ,
         \CARRYB[11][14] , \CARRYB[11][13] , \CARRYB[11][12] ,
         \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] , \CARRYB[11][8] ,
         \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[11][0] ,
         \CARRYB[10][14] , \CARRYB[10][13] , \CARRYB[10][12] ,
         \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] ,
         \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] , \CARRYB[10][4] ,
         \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] , \CARRYB[10][0] ,
         \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] , \CARRYB[9][11] ,
         \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] , \CARRYB[9][7] ,
         \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] , \CARRYB[8][14] ,
         \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] ,
         \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] ,
         \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] ,
         \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] ,
         \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] ,
         \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] , \CARRYB[6][4] ,
         \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] , \CARRYB[6][0] ,
         \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] ,
         \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] ,
         \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][14] ,
         \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] ,
         \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][6] ,
         \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] , \CARRYB[4][2] ,
         \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][14] , \CARRYB[3][13] ,
         \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] , \CARRYB[3][9] ,
         \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[3][0] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[15][0] , \SUMB[14][14] ,
         \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] ,
         \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] ,
         \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] ,
         \SUMB[14][1] , \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] ,
         \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] ,
         \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] ,
         \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][14] ,
         \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] ,
         \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] ,
         \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] ,
         \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] ,
         \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] ,
         \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] ,
         \SUMB[10][1] , \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] ,
         \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] ,
         \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] ,
         \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] , \SUMB[8][13] ,
         \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] , \SUMB[8][9] ,
         \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] , \SUMB[6][5] ,
         \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] ,
         \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] , \SUMB[4][5] ,
         \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] ,
         \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] , \A1[28] ,
         \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] ,
         \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] ,
         \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] ,
         \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64;
  wire   SYNOPSYS_UNCONNECTED__0;

  FADDX1 S4_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), .CO(
        \CARRYB[15][0] ), .S(\SUMB[15][0] ) );
  FADDX1 S4_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FADDX1 S4_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FADDX1 S4_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FADDX1 S4_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1 S4_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), .CO(
        \CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FADDX1 S4_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FADDX1 S4_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FADDX1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FADDX1 S4_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FADDX1 S4_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FADDX1 S4_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1 S4_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1 S5_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\ab[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FADDX1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FADDX1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FADDX1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FADDX1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FADDX1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FADDX1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FADDX1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FADDX1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FADDX1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FADDX1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1 S3_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\ab[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FADDX1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FADDX1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FADDX1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FADDX1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FADDX1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FADDX1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FADDX1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FADDX1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FADDX1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FADDX1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FADDX1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FADDX1 S3_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\ab[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FADDX1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FADDX1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FADDX1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FADDX1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FADDX1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FADDX1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FADDX1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FADDX1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FADDX1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FADDX1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FADDX1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FADDX1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FADDX1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FADDX1 S3_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\ab[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FADDX1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FADDX1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FADDX1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FADDX1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FADDX1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FADDX1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FADDX1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FADDX1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FADDX1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FADDX1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FADDX1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FADDX1 S3_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\ab[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FADDX1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), 
        .CO(\CARRYB[10][0] ), .S(\A1[8] ) );
  FADDX1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), 
        .CO(\CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FADDX1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), 
        .CO(\CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FADDX1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), 
        .CO(\CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FADDX1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), 
        .CO(\CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FADDX1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), 
        .CO(\CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FADDX1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FADDX1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FADDX1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FADDX1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FADDX1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FADDX1 S3_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\ab[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FADDX1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FADDX1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FADDX1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FADDX1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FADDX1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FADDX1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FADDX1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FADDX1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FADDX1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FADDX1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FADDX1 S3_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\ab[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FADDX1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FADDX1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FADDX1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FADDX1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FADDX1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FADDX1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FADDX1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FADDX1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FADDX1 S3_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\ab[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FADDX1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FADDX1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FADDX1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FADDX1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FADDX1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FADDX1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FADDX1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FADDX1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FADDX1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FADDX1 S3_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\ab[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FADDX1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FADDX1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FADDX1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FADDX1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FADDX1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FADDX1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FADDX1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FADDX1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FADDX1 S3_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\ab[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FADDX1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FADDX1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FADDX1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FADDX1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FADDX1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FADDX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FADDX1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FADDX1 S3_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\ab[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FADDX1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FADDX1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FADDX1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FADDX1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FADDX1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FADDX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FADDX1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FADDX1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FADDX1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FADDX1 S3_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\ab[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FADDX1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FADDX1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FADDX1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FADDX1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FADDX1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FADDX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FADDX1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FADDX1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FADDX1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FADDX1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1 S3_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\ab[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FADDX1 S1_2_0 ( .A(\ab[2][0] ), .B(n18), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FADDX1 S2_2_1 ( .A(\ab[2][1] ), .B(n17), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1 S2_2_2 ( .A(\ab[2][2] ), .B(n16), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FADDX1 S2_2_3 ( .A(\ab[2][3] ), .B(n15), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1 S2_2_4 ( .A(\ab[2][4] ), .B(n14), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1 S2_2_5 ( .A(\ab[2][5] ), .B(n13), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FADDX1 S2_2_6 ( .A(\ab[2][6] ), .B(n12), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FADDX1 S2_2_7 ( .A(\ab[2][7] ), .B(n11), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FADDX1 S2_2_8 ( .A(\ab[2][8] ), .B(n10), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FADDX1 S2_2_9 ( .A(\ab[2][9] ), .B(n9), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1 S2_2_10 ( .A(\ab[2][10] ), .B(n8), .CI(\SUMB[1][11] ), .CO(
        \CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FADDX1 S2_2_11 ( .A(\ab[2][11] ), .B(n7), .CI(\SUMB[1][12] ), .CO(
        \CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1 S2_2_12 ( .A(\ab[2][12] ), .B(n6), .CI(\SUMB[1][13] ), .CO(
        \CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FADDX1 S2_2_13 ( .A(\ab[2][13] ), .B(n5), .CI(\SUMB[1][14] ), .CO(
        \CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FADDX1 S3_2_14 ( .A(\ab[2][14] ), .B(n4), .CI(\ab[1][15] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  betterNeighborsInMyCluster_DW01_add_10 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , 
        \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , 
        \SUMB[15][0] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , 
        \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({
        n3, n19, n27, n32, n26, n25, n30, n31, n29, n28, n24, n23, n21, n22, 
        n20, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        PRODUCT[30:2]}) );
  AND2X1 U2 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[15][15] ), .Q(n3) );
  AND2X1 U3 ( .IN1(\ab[0][15] ), .IN2(\ab[1][14] ), .Q(n4) );
  AND2X1 U4 ( .IN1(\ab[0][14] ), .IN2(\ab[1][13] ), .Q(n5) );
  AND2X1 U5 ( .IN1(\ab[0][13] ), .IN2(\ab[1][12] ), .Q(n6) );
  AND2X1 U6 ( .IN1(\ab[0][12] ), .IN2(\ab[1][11] ), .Q(n7) );
  AND2X1 U7 ( .IN1(\ab[0][11] ), .IN2(\ab[1][10] ), .Q(n8) );
  AND2X1 U8 ( .IN1(\ab[0][10] ), .IN2(\ab[1][9] ), .Q(n9) );
  AND2X1 U9 ( .IN1(\ab[0][9] ), .IN2(\ab[1][8] ), .Q(n10) );
  AND2X1 U10 ( .IN1(\ab[0][8] ), .IN2(\ab[1][7] ), .Q(n11) );
  AND2X1 U11 ( .IN1(\ab[0][7] ), .IN2(\ab[1][6] ), .Q(n12) );
  AND2X1 U12 ( .IN1(\ab[0][6] ), .IN2(\ab[1][5] ), .Q(n13) );
  AND2X1 U13 ( .IN1(\ab[0][5] ), .IN2(\ab[1][4] ), .Q(n14) );
  AND2X1 U14 ( .IN1(\ab[0][4] ), .IN2(\ab[1][3] ), .Q(n15) );
  AND2X1 U15 ( .IN1(\ab[0][3] ), .IN2(\ab[1][2] ), .Q(n16) );
  AND2X1 U16 ( .IN1(\ab[0][2] ), .IN2(\ab[1][1] ), .Q(n17) );
  AND2X1 U17 ( .IN1(\ab[0][1] ), .IN2(\ab[1][0] ), .Q(n18) );
  AND2X1 U18 ( .IN1(\CARRYB[15][13] ), .IN2(\SUMB[15][14] ), .Q(n19) );
  AND2X1 U19 ( .IN1(\CARRYB[15][0] ), .IN2(\SUMB[15][1] ), .Q(n20) );
  AND2X1 U20 ( .IN1(\CARRYB[15][2] ), .IN2(\SUMB[15][3] ), .Q(n21) );
  AND2X1 U21 ( .IN1(\CARRYB[15][1] ), .IN2(\SUMB[15][2] ), .Q(n22) );
  AND2X1 U22 ( .IN1(\CARRYB[15][3] ), .IN2(\SUMB[15][4] ), .Q(n23) );
  AND2X1 U23 ( .IN1(\CARRYB[15][4] ), .IN2(\SUMB[15][5] ), .Q(n24) );
  AND2X1 U24 ( .IN1(\CARRYB[15][9] ), .IN2(\SUMB[15][10] ), .Q(n25) );
  AND2X1 U25 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .Q(n26) );
  AND2X1 U26 ( .IN1(\CARRYB[15][12] ), .IN2(\SUMB[15][13] ), .Q(n27) );
  AND2X1 U27 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[15][6] ), .Q(n28) );
  AND2X1 U28 ( .IN1(\CARRYB[15][6] ), .IN2(\SUMB[15][7] ), .Q(n29) );
  AND2X1 U29 ( .IN1(\CARRYB[15][8] ), .IN2(\SUMB[15][9] ), .Q(n30) );
  AND2X1 U30 ( .IN1(\CARRYB[15][7] ), .IN2(\SUMB[15][8] ), .Q(n31) );
  AND2X1 U31 ( .IN1(\CARRYB[15][11] ), .IN2(\SUMB[15][12] ), .Q(n32) );
  INVX0 U32 ( .INP(B[7]), .ZN(n41) );
  INVX0 U33 ( .INP(B[1]), .ZN(n47) );
  INVX0 U34 ( .INP(B[2]), .ZN(n46) );
  INVX0 U35 ( .INP(B[3]), .ZN(n45) );
  INVX0 U36 ( .INP(B[6]), .ZN(n42) );
  INVX0 U37 ( .INP(B[8]), .ZN(n40) );
  INVX0 U38 ( .INP(B[9]), .ZN(n39) );
  INVX0 U39 ( .INP(B[10]), .ZN(n38) );
  INVX0 U40 ( .INP(B[11]), .ZN(n37) );
  INVX0 U41 ( .INP(B[5]), .ZN(n43) );
  INVX0 U42 ( .INP(B[4]), .ZN(n44) );
  INVX0 U43 ( .INP(B[0]), .ZN(n48) );
  INVX0 U44 ( .INP(B[12]), .ZN(n36) );
  INVX0 U45 ( .INP(B[13]), .ZN(n35) );
  INVX0 U46 ( .INP(B[14]), .ZN(n34) );
  INVX0 U47 ( .INP(B[15]), .ZN(n33) );
  INVX0 U48 ( .INP(A[0]), .ZN(n64) );
  INVX0 U49 ( .INP(A[3]), .ZN(n61) );
  INVX0 U50 ( .INP(A[1]), .ZN(n63) );
  INVX0 U51 ( .INP(A[4]), .ZN(n60) );
  INVX0 U52 ( .INP(A[5]), .ZN(n59) );
  INVX0 U53 ( .INP(A[2]), .ZN(n62) );
  INVX0 U54 ( .INP(A[6]), .ZN(n58) );
  INVX0 U55 ( .INP(A[9]), .ZN(n55) );
  INVX0 U56 ( .INP(A[7]), .ZN(n57) );
  INVX0 U57 ( .INP(A[8]), .ZN(n56) );
  INVX0 U58 ( .INP(A[10]), .ZN(n54) );
  INVX0 U59 ( .INP(A[11]), .ZN(n53) );
  INVX0 U60 ( .INP(A[12]), .ZN(n52) );
  INVX0 U61 ( .INP(A[13]), .ZN(n51) );
  INVX0 U62 ( .INP(A[14]), .ZN(n50) );
  INVX0 U63 ( .INP(A[15]), .ZN(n49) );
  XOR2X1 U64 ( .IN1(\CARRYB[15][0] ), .IN2(\SUMB[15][1] ), .Q(\A1[14] ) );
  XOR2X1 U65 ( .IN1(\CARRYB[15][1] ), .IN2(\SUMB[15][2] ), .Q(\A1[15] ) );
  XOR2X1 U66 ( .IN1(\CARRYB[15][2] ), .IN2(\SUMB[15][3] ), .Q(\A1[16] ) );
  XOR2X1 U67 ( .IN1(\CARRYB[15][3] ), .IN2(\SUMB[15][4] ), .Q(\A1[17] ) );
  XOR2X1 U68 ( .IN1(\CARRYB[15][4] ), .IN2(\SUMB[15][5] ), .Q(\A1[18] ) );
  XOR2X1 U69 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[15][6] ), .Q(\A1[19] ) );
  XOR2X1 U70 ( .IN1(\CARRYB[15][6] ), .IN2(\SUMB[15][7] ), .Q(\A1[20] ) );
  XOR2X1 U71 ( .IN1(\CARRYB[15][7] ), .IN2(\SUMB[15][8] ), .Q(\A1[21] ) );
  XOR2X1 U72 ( .IN1(\CARRYB[15][8] ), .IN2(\SUMB[15][9] ), .Q(\A1[22] ) );
  XOR2X1 U73 ( .IN1(\CARRYB[15][9] ), .IN2(\SUMB[15][10] ), .Q(\A1[23] ) );
  XOR2X1 U74 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .Q(\A1[24] ) );
  XOR2X1 U75 ( .IN1(\CARRYB[15][11] ), .IN2(\SUMB[15][12] ), .Q(\A1[25] ) );
  XOR2X1 U76 ( .IN1(\CARRYB[15][12] ), .IN2(\SUMB[15][13] ), .Q(\A1[26] ) );
  XOR2X1 U77 ( .IN1(\CARRYB[15][13] ), .IN2(\SUMB[15][14] ), .Q(\A1[27] ) );
  XOR2X1 U78 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[15][15] ), .Q(\A1[28] ) );
  XOR2X1 U79 ( .IN1(\ab[1][0] ), .IN2(\ab[0][1] ), .Q(PRODUCT[1]) );
  XOR2X1 U80 ( .IN1(\ab[1][1] ), .IN2(\ab[0][2] ), .Q(\SUMB[1][1] ) );
  XOR2X1 U81 ( .IN1(\ab[1][2] ), .IN2(\ab[0][3] ), .Q(\SUMB[1][2] ) );
  XOR2X1 U82 ( .IN1(\ab[1][3] ), .IN2(\ab[0][4] ), .Q(\SUMB[1][3] ) );
  XOR2X1 U83 ( .IN1(\ab[1][4] ), .IN2(\ab[0][5] ), .Q(\SUMB[1][4] ) );
  XOR2X1 U84 ( .IN1(\ab[1][5] ), .IN2(\ab[0][6] ), .Q(\SUMB[1][5] ) );
  XOR2X1 U85 ( .IN1(\ab[1][6] ), .IN2(\ab[0][7] ), .Q(\SUMB[1][6] ) );
  XOR2X1 U86 ( .IN1(\ab[1][7] ), .IN2(\ab[0][8] ), .Q(\SUMB[1][7] ) );
  XOR2X1 U87 ( .IN1(\ab[1][8] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][8] ) );
  XOR2X1 U88 ( .IN1(\ab[1][9] ), .IN2(\ab[0][10] ), .Q(\SUMB[1][9] ) );
  XOR2X1 U89 ( .IN1(\ab[1][10] ), .IN2(\ab[0][11] ), .Q(\SUMB[1][10] ) );
  XOR2X1 U90 ( .IN1(\ab[1][11] ), .IN2(\ab[0][12] ), .Q(\SUMB[1][11] ) );
  XOR2X1 U91 ( .IN1(\ab[1][12] ), .IN2(\ab[0][13] ), .Q(\SUMB[1][12] ) );
  XOR2X1 U92 ( .IN1(\ab[1][13] ), .IN2(\ab[0][14] ), .Q(\SUMB[1][13] ) );
  XOR2X1 U93 ( .IN1(\ab[1][14] ), .IN2(\ab[0][15] ), .Q(\SUMB[1][14] ) );
  NOR2X0 U95 ( .IN1(n55), .IN2(n39), .QN(\ab[9][9] ) );
  NOR2X0 U96 ( .IN1(n55), .IN2(n40), .QN(\ab[9][8] ) );
  NOR2X0 U97 ( .IN1(n55), .IN2(n41), .QN(\ab[9][7] ) );
  NOR2X0 U98 ( .IN1(n55), .IN2(n42), .QN(\ab[9][6] ) );
  NOR2X0 U99 ( .IN1(n55), .IN2(n43), .QN(\ab[9][5] ) );
  NOR2X0 U100 ( .IN1(n55), .IN2(n44), .QN(\ab[9][4] ) );
  NOR2X0 U101 ( .IN1(n55), .IN2(n45), .QN(\ab[9][3] ) );
  NOR2X0 U102 ( .IN1(n55), .IN2(n46), .QN(\ab[9][2] ) );
  NOR2X0 U103 ( .IN1(n55), .IN2(n47), .QN(\ab[9][1] ) );
  NOR2X0 U104 ( .IN1(n55), .IN2(n33), .QN(\ab[9][15] ) );
  NOR2X0 U105 ( .IN1(n55), .IN2(n34), .QN(\ab[9][14] ) );
  NOR2X0 U106 ( .IN1(n55), .IN2(n35), .QN(\ab[9][13] ) );
  NOR2X0 U107 ( .IN1(n55), .IN2(n36), .QN(\ab[9][12] ) );
  NOR2X0 U108 ( .IN1(n55), .IN2(n37), .QN(\ab[9][11] ) );
  NOR2X0 U109 ( .IN1(n55), .IN2(n38), .QN(\ab[9][10] ) );
  NOR2X0 U110 ( .IN1(n55), .IN2(n48), .QN(\ab[9][0] ) );
  NOR2X0 U111 ( .IN1(n39), .IN2(n56), .QN(\ab[8][9] ) );
  NOR2X0 U112 ( .IN1(n40), .IN2(n56), .QN(\ab[8][8] ) );
  NOR2X0 U113 ( .IN1(n41), .IN2(n56), .QN(\ab[8][7] ) );
  NOR2X0 U114 ( .IN1(n42), .IN2(n56), .QN(\ab[8][6] ) );
  NOR2X0 U115 ( .IN1(n43), .IN2(n56), .QN(\ab[8][5] ) );
  NOR2X0 U116 ( .IN1(n44), .IN2(n56), .QN(\ab[8][4] ) );
  NOR2X0 U117 ( .IN1(n45), .IN2(n56), .QN(\ab[8][3] ) );
  NOR2X0 U118 ( .IN1(n46), .IN2(n56), .QN(\ab[8][2] ) );
  NOR2X0 U119 ( .IN1(n47), .IN2(n56), .QN(\ab[8][1] ) );
  NOR2X0 U120 ( .IN1(n33), .IN2(n56), .QN(\ab[8][15] ) );
  NOR2X0 U121 ( .IN1(n34), .IN2(n56), .QN(\ab[8][14] ) );
  NOR2X0 U122 ( .IN1(n35), .IN2(n56), .QN(\ab[8][13] ) );
  NOR2X0 U123 ( .IN1(n36), .IN2(n56), .QN(\ab[8][12] ) );
  NOR2X0 U124 ( .IN1(n37), .IN2(n56), .QN(\ab[8][11] ) );
  NOR2X0 U125 ( .IN1(n38), .IN2(n56), .QN(\ab[8][10] ) );
  NOR2X0 U126 ( .IN1(n48), .IN2(n56), .QN(\ab[8][0] ) );
  NOR2X0 U127 ( .IN1(n39), .IN2(n57), .QN(\ab[7][9] ) );
  NOR2X0 U128 ( .IN1(n40), .IN2(n57), .QN(\ab[7][8] ) );
  NOR2X0 U129 ( .IN1(n41), .IN2(n57), .QN(\ab[7][7] ) );
  NOR2X0 U130 ( .IN1(n42), .IN2(n57), .QN(\ab[7][6] ) );
  NOR2X0 U131 ( .IN1(n43), .IN2(n57), .QN(\ab[7][5] ) );
  NOR2X0 U132 ( .IN1(n44), .IN2(n57), .QN(\ab[7][4] ) );
  NOR2X0 U133 ( .IN1(n45), .IN2(n57), .QN(\ab[7][3] ) );
  NOR2X0 U134 ( .IN1(n46), .IN2(n57), .QN(\ab[7][2] ) );
  NOR2X0 U135 ( .IN1(n47), .IN2(n57), .QN(\ab[7][1] ) );
  NOR2X0 U136 ( .IN1(n33), .IN2(n57), .QN(\ab[7][15] ) );
  NOR2X0 U137 ( .IN1(n34), .IN2(n57), .QN(\ab[7][14] ) );
  NOR2X0 U138 ( .IN1(n35), .IN2(n57), .QN(\ab[7][13] ) );
  NOR2X0 U139 ( .IN1(n36), .IN2(n57), .QN(\ab[7][12] ) );
  NOR2X0 U140 ( .IN1(n37), .IN2(n57), .QN(\ab[7][11] ) );
  NOR2X0 U141 ( .IN1(n38), .IN2(n57), .QN(\ab[7][10] ) );
  NOR2X0 U142 ( .IN1(n48), .IN2(n57), .QN(\ab[7][0] ) );
  NOR2X0 U143 ( .IN1(n39), .IN2(n58), .QN(\ab[6][9] ) );
  NOR2X0 U144 ( .IN1(n40), .IN2(n58), .QN(\ab[6][8] ) );
  NOR2X0 U145 ( .IN1(n41), .IN2(n58), .QN(\ab[6][7] ) );
  NOR2X0 U146 ( .IN1(n42), .IN2(n58), .QN(\ab[6][6] ) );
  NOR2X0 U147 ( .IN1(n43), .IN2(n58), .QN(\ab[6][5] ) );
  NOR2X0 U148 ( .IN1(n44), .IN2(n58), .QN(\ab[6][4] ) );
  NOR2X0 U149 ( .IN1(n45), .IN2(n58), .QN(\ab[6][3] ) );
  NOR2X0 U150 ( .IN1(n46), .IN2(n58), .QN(\ab[6][2] ) );
  NOR2X0 U151 ( .IN1(n47), .IN2(n58), .QN(\ab[6][1] ) );
  NOR2X0 U152 ( .IN1(n33), .IN2(n58), .QN(\ab[6][15] ) );
  NOR2X0 U153 ( .IN1(n34), .IN2(n58), .QN(\ab[6][14] ) );
  NOR2X0 U154 ( .IN1(n35), .IN2(n58), .QN(\ab[6][13] ) );
  NOR2X0 U155 ( .IN1(n36), .IN2(n58), .QN(\ab[6][12] ) );
  NOR2X0 U156 ( .IN1(n37), .IN2(n58), .QN(\ab[6][11] ) );
  NOR2X0 U157 ( .IN1(n38), .IN2(n58), .QN(\ab[6][10] ) );
  NOR2X0 U158 ( .IN1(n48), .IN2(n58), .QN(\ab[6][0] ) );
  NOR2X0 U159 ( .IN1(n39), .IN2(n59), .QN(\ab[5][9] ) );
  NOR2X0 U160 ( .IN1(n40), .IN2(n59), .QN(\ab[5][8] ) );
  NOR2X0 U161 ( .IN1(n41), .IN2(n59), .QN(\ab[5][7] ) );
  NOR2X0 U162 ( .IN1(n42), .IN2(n59), .QN(\ab[5][6] ) );
  NOR2X0 U163 ( .IN1(n43), .IN2(n59), .QN(\ab[5][5] ) );
  NOR2X0 U164 ( .IN1(n44), .IN2(n59), .QN(\ab[5][4] ) );
  NOR2X0 U165 ( .IN1(n45), .IN2(n59), .QN(\ab[5][3] ) );
  NOR2X0 U166 ( .IN1(n46), .IN2(n59), .QN(\ab[5][2] ) );
  NOR2X0 U167 ( .IN1(n47), .IN2(n59), .QN(\ab[5][1] ) );
  NOR2X0 U168 ( .IN1(n33), .IN2(n59), .QN(\ab[5][15] ) );
  NOR2X0 U169 ( .IN1(n34), .IN2(n59), .QN(\ab[5][14] ) );
  NOR2X0 U170 ( .IN1(n35), .IN2(n59), .QN(\ab[5][13] ) );
  NOR2X0 U171 ( .IN1(n36), .IN2(n59), .QN(\ab[5][12] ) );
  NOR2X0 U172 ( .IN1(n37), .IN2(n59), .QN(\ab[5][11] ) );
  NOR2X0 U173 ( .IN1(n38), .IN2(n59), .QN(\ab[5][10] ) );
  NOR2X0 U174 ( .IN1(n48), .IN2(n59), .QN(\ab[5][0] ) );
  NOR2X0 U175 ( .IN1(n39), .IN2(n60), .QN(\ab[4][9] ) );
  NOR2X0 U176 ( .IN1(n40), .IN2(n60), .QN(\ab[4][8] ) );
  NOR2X0 U177 ( .IN1(n41), .IN2(n60), .QN(\ab[4][7] ) );
  NOR2X0 U178 ( .IN1(n42), .IN2(n60), .QN(\ab[4][6] ) );
  NOR2X0 U179 ( .IN1(n43), .IN2(n60), .QN(\ab[4][5] ) );
  NOR2X0 U180 ( .IN1(n44), .IN2(n60), .QN(\ab[4][4] ) );
  NOR2X0 U181 ( .IN1(n45), .IN2(n60), .QN(\ab[4][3] ) );
  NOR2X0 U182 ( .IN1(n46), .IN2(n60), .QN(\ab[4][2] ) );
  NOR2X0 U183 ( .IN1(n47), .IN2(n60), .QN(\ab[4][1] ) );
  NOR2X0 U184 ( .IN1(n33), .IN2(n60), .QN(\ab[4][15] ) );
  NOR2X0 U185 ( .IN1(n34), .IN2(n60), .QN(\ab[4][14] ) );
  NOR2X0 U186 ( .IN1(n35), .IN2(n60), .QN(\ab[4][13] ) );
  NOR2X0 U187 ( .IN1(n36), .IN2(n60), .QN(\ab[4][12] ) );
  NOR2X0 U188 ( .IN1(n37), .IN2(n60), .QN(\ab[4][11] ) );
  NOR2X0 U189 ( .IN1(n38), .IN2(n60), .QN(\ab[4][10] ) );
  NOR2X0 U190 ( .IN1(n48), .IN2(n60), .QN(\ab[4][0] ) );
  NOR2X0 U191 ( .IN1(n39), .IN2(n61), .QN(\ab[3][9] ) );
  NOR2X0 U192 ( .IN1(n40), .IN2(n61), .QN(\ab[3][8] ) );
  NOR2X0 U193 ( .IN1(n41), .IN2(n61), .QN(\ab[3][7] ) );
  NOR2X0 U194 ( .IN1(n42), .IN2(n61), .QN(\ab[3][6] ) );
  NOR2X0 U195 ( .IN1(n43), .IN2(n61), .QN(\ab[3][5] ) );
  NOR2X0 U196 ( .IN1(n44), .IN2(n61), .QN(\ab[3][4] ) );
  NOR2X0 U197 ( .IN1(n45), .IN2(n61), .QN(\ab[3][3] ) );
  NOR2X0 U198 ( .IN1(n46), .IN2(n61), .QN(\ab[3][2] ) );
  NOR2X0 U199 ( .IN1(n47), .IN2(n61), .QN(\ab[3][1] ) );
  NOR2X0 U200 ( .IN1(n33), .IN2(n61), .QN(\ab[3][15] ) );
  NOR2X0 U201 ( .IN1(n34), .IN2(n61), .QN(\ab[3][14] ) );
  NOR2X0 U202 ( .IN1(n35), .IN2(n61), .QN(\ab[3][13] ) );
  NOR2X0 U203 ( .IN1(n36), .IN2(n61), .QN(\ab[3][12] ) );
  NOR2X0 U204 ( .IN1(n37), .IN2(n61), .QN(\ab[3][11] ) );
  NOR2X0 U205 ( .IN1(n38), .IN2(n61), .QN(\ab[3][10] ) );
  NOR2X0 U206 ( .IN1(n48), .IN2(n61), .QN(\ab[3][0] ) );
  NOR2X0 U207 ( .IN1(n39), .IN2(n62), .QN(\ab[2][9] ) );
  NOR2X0 U208 ( .IN1(n40), .IN2(n62), .QN(\ab[2][8] ) );
  NOR2X0 U209 ( .IN1(n41), .IN2(n62), .QN(\ab[2][7] ) );
  NOR2X0 U210 ( .IN1(n42), .IN2(n62), .QN(\ab[2][6] ) );
  NOR2X0 U211 ( .IN1(n43), .IN2(n62), .QN(\ab[2][5] ) );
  NOR2X0 U212 ( .IN1(n44), .IN2(n62), .QN(\ab[2][4] ) );
  NOR2X0 U213 ( .IN1(n45), .IN2(n62), .QN(\ab[2][3] ) );
  NOR2X0 U214 ( .IN1(n46), .IN2(n62), .QN(\ab[2][2] ) );
  NOR2X0 U215 ( .IN1(n47), .IN2(n62), .QN(\ab[2][1] ) );
  NOR2X0 U216 ( .IN1(n33), .IN2(n62), .QN(\ab[2][15] ) );
  NOR2X0 U217 ( .IN1(n34), .IN2(n62), .QN(\ab[2][14] ) );
  NOR2X0 U218 ( .IN1(n35), .IN2(n62), .QN(\ab[2][13] ) );
  NOR2X0 U219 ( .IN1(n36), .IN2(n62), .QN(\ab[2][12] ) );
  NOR2X0 U220 ( .IN1(n37), .IN2(n62), .QN(\ab[2][11] ) );
  NOR2X0 U221 ( .IN1(n38), .IN2(n62), .QN(\ab[2][10] ) );
  NOR2X0 U222 ( .IN1(n48), .IN2(n62), .QN(\ab[2][0] ) );
  NOR2X0 U223 ( .IN1(n39), .IN2(n63), .QN(\ab[1][9] ) );
  NOR2X0 U224 ( .IN1(n40), .IN2(n63), .QN(\ab[1][8] ) );
  NOR2X0 U225 ( .IN1(n41), .IN2(n63), .QN(\ab[1][7] ) );
  NOR2X0 U226 ( .IN1(n42), .IN2(n63), .QN(\ab[1][6] ) );
  NOR2X0 U227 ( .IN1(n43), .IN2(n63), .QN(\ab[1][5] ) );
  NOR2X0 U228 ( .IN1(n44), .IN2(n63), .QN(\ab[1][4] ) );
  NOR2X0 U229 ( .IN1(n45), .IN2(n63), .QN(\ab[1][3] ) );
  NOR2X0 U230 ( .IN1(n46), .IN2(n63), .QN(\ab[1][2] ) );
  NOR2X0 U231 ( .IN1(n47), .IN2(n63), .QN(\ab[1][1] ) );
  NOR2X0 U232 ( .IN1(n33), .IN2(n63), .QN(\ab[1][15] ) );
  NOR2X0 U233 ( .IN1(n34), .IN2(n63), .QN(\ab[1][14] ) );
  NOR2X0 U234 ( .IN1(n35), .IN2(n63), .QN(\ab[1][13] ) );
  NOR2X0 U235 ( .IN1(n36), .IN2(n63), .QN(\ab[1][12] ) );
  NOR2X0 U236 ( .IN1(n37), .IN2(n63), .QN(\ab[1][11] ) );
  NOR2X0 U237 ( .IN1(n38), .IN2(n63), .QN(\ab[1][10] ) );
  NOR2X0 U238 ( .IN1(n48), .IN2(n63), .QN(\ab[1][0] ) );
  NOR2X0 U239 ( .IN1(n39), .IN2(n49), .QN(\ab[15][9] ) );
  NOR2X0 U240 ( .IN1(n40), .IN2(n49), .QN(\ab[15][8] ) );
  NOR2X0 U241 ( .IN1(n41), .IN2(n49), .QN(\ab[15][7] ) );
  NOR2X0 U242 ( .IN1(n42), .IN2(n49), .QN(\ab[15][6] ) );
  NOR2X0 U243 ( .IN1(n43), .IN2(n49), .QN(\ab[15][5] ) );
  NOR2X0 U244 ( .IN1(n44), .IN2(n49), .QN(\ab[15][4] ) );
  NOR2X0 U245 ( .IN1(n45), .IN2(n49), .QN(\ab[15][3] ) );
  NOR2X0 U246 ( .IN1(n46), .IN2(n49), .QN(\ab[15][2] ) );
  NOR2X0 U247 ( .IN1(n47), .IN2(n49), .QN(\ab[15][1] ) );
  NOR2X0 U248 ( .IN1(n33), .IN2(n49), .QN(\ab[15][15] ) );
  NOR2X0 U249 ( .IN1(n34), .IN2(n49), .QN(\ab[15][14] ) );
  NOR2X0 U250 ( .IN1(n35), .IN2(n49), .QN(\ab[15][13] ) );
  NOR2X0 U251 ( .IN1(n36), .IN2(n49), .QN(\ab[15][12] ) );
  NOR2X0 U252 ( .IN1(n37), .IN2(n49), .QN(\ab[15][11] ) );
  NOR2X0 U253 ( .IN1(n38), .IN2(n49), .QN(\ab[15][10] ) );
  NOR2X0 U254 ( .IN1(n48), .IN2(n49), .QN(\ab[15][0] ) );
  NOR2X0 U255 ( .IN1(n39), .IN2(n50), .QN(\ab[14][9] ) );
  NOR2X0 U256 ( .IN1(n40), .IN2(n50), .QN(\ab[14][8] ) );
  NOR2X0 U257 ( .IN1(n41), .IN2(n50), .QN(\ab[14][7] ) );
  NOR2X0 U258 ( .IN1(n42), .IN2(n50), .QN(\ab[14][6] ) );
  NOR2X0 U259 ( .IN1(n43), .IN2(n50), .QN(\ab[14][5] ) );
  NOR2X0 U260 ( .IN1(n44), .IN2(n50), .QN(\ab[14][4] ) );
  NOR2X0 U261 ( .IN1(n45), .IN2(n50), .QN(\ab[14][3] ) );
  NOR2X0 U262 ( .IN1(n46), .IN2(n50), .QN(\ab[14][2] ) );
  NOR2X0 U263 ( .IN1(n47), .IN2(n50), .QN(\ab[14][1] ) );
  NOR2X0 U264 ( .IN1(n33), .IN2(n50), .QN(\ab[14][15] ) );
  NOR2X0 U265 ( .IN1(n34), .IN2(n50), .QN(\ab[14][14] ) );
  NOR2X0 U266 ( .IN1(n35), .IN2(n50), .QN(\ab[14][13] ) );
  NOR2X0 U267 ( .IN1(n36), .IN2(n50), .QN(\ab[14][12] ) );
  NOR2X0 U268 ( .IN1(n37), .IN2(n50), .QN(\ab[14][11] ) );
  NOR2X0 U269 ( .IN1(n38), .IN2(n50), .QN(\ab[14][10] ) );
  NOR2X0 U270 ( .IN1(n48), .IN2(n50), .QN(\ab[14][0] ) );
  NOR2X0 U271 ( .IN1(n39), .IN2(n51), .QN(\ab[13][9] ) );
  NOR2X0 U272 ( .IN1(n40), .IN2(n51), .QN(\ab[13][8] ) );
  NOR2X0 U273 ( .IN1(n41), .IN2(n51), .QN(\ab[13][7] ) );
  NOR2X0 U274 ( .IN1(n42), .IN2(n51), .QN(\ab[13][6] ) );
  NOR2X0 U275 ( .IN1(n43), .IN2(n51), .QN(\ab[13][5] ) );
  NOR2X0 U276 ( .IN1(n44), .IN2(n51), .QN(\ab[13][4] ) );
  NOR2X0 U277 ( .IN1(n45), .IN2(n51), .QN(\ab[13][3] ) );
  NOR2X0 U278 ( .IN1(n46), .IN2(n51), .QN(\ab[13][2] ) );
  NOR2X0 U279 ( .IN1(n47), .IN2(n51), .QN(\ab[13][1] ) );
  NOR2X0 U280 ( .IN1(n33), .IN2(n51), .QN(\ab[13][15] ) );
  NOR2X0 U281 ( .IN1(n34), .IN2(n51), .QN(\ab[13][14] ) );
  NOR2X0 U282 ( .IN1(n35), .IN2(n51), .QN(\ab[13][13] ) );
  NOR2X0 U283 ( .IN1(n36), .IN2(n51), .QN(\ab[13][12] ) );
  NOR2X0 U284 ( .IN1(n37), .IN2(n51), .QN(\ab[13][11] ) );
  NOR2X0 U285 ( .IN1(n38), .IN2(n51), .QN(\ab[13][10] ) );
  NOR2X0 U286 ( .IN1(n48), .IN2(n51), .QN(\ab[13][0] ) );
  NOR2X0 U287 ( .IN1(n39), .IN2(n52), .QN(\ab[12][9] ) );
  NOR2X0 U288 ( .IN1(n40), .IN2(n52), .QN(\ab[12][8] ) );
  NOR2X0 U289 ( .IN1(n41), .IN2(n52), .QN(\ab[12][7] ) );
  NOR2X0 U290 ( .IN1(n42), .IN2(n52), .QN(\ab[12][6] ) );
  NOR2X0 U291 ( .IN1(n43), .IN2(n52), .QN(\ab[12][5] ) );
  NOR2X0 U292 ( .IN1(n44), .IN2(n52), .QN(\ab[12][4] ) );
  NOR2X0 U293 ( .IN1(n45), .IN2(n52), .QN(\ab[12][3] ) );
  NOR2X0 U294 ( .IN1(n46), .IN2(n52), .QN(\ab[12][2] ) );
  NOR2X0 U295 ( .IN1(n47), .IN2(n52), .QN(\ab[12][1] ) );
  NOR2X0 U296 ( .IN1(n33), .IN2(n52), .QN(\ab[12][15] ) );
  NOR2X0 U297 ( .IN1(n34), .IN2(n52), .QN(\ab[12][14] ) );
  NOR2X0 U298 ( .IN1(n35), .IN2(n52), .QN(\ab[12][13] ) );
  NOR2X0 U299 ( .IN1(n36), .IN2(n52), .QN(\ab[12][12] ) );
  NOR2X0 U300 ( .IN1(n37), .IN2(n52), .QN(\ab[12][11] ) );
  NOR2X0 U301 ( .IN1(n38), .IN2(n52), .QN(\ab[12][10] ) );
  NOR2X0 U302 ( .IN1(n48), .IN2(n52), .QN(\ab[12][0] ) );
  NOR2X0 U303 ( .IN1(n39), .IN2(n53), .QN(\ab[11][9] ) );
  NOR2X0 U304 ( .IN1(n40), .IN2(n53), .QN(\ab[11][8] ) );
  NOR2X0 U305 ( .IN1(n41), .IN2(n53), .QN(\ab[11][7] ) );
  NOR2X0 U306 ( .IN1(n42), .IN2(n53), .QN(\ab[11][6] ) );
  NOR2X0 U307 ( .IN1(n43), .IN2(n53), .QN(\ab[11][5] ) );
  NOR2X0 U308 ( .IN1(n44), .IN2(n53), .QN(\ab[11][4] ) );
  NOR2X0 U309 ( .IN1(n45), .IN2(n53), .QN(\ab[11][3] ) );
  NOR2X0 U310 ( .IN1(n46), .IN2(n53), .QN(\ab[11][2] ) );
  NOR2X0 U311 ( .IN1(n47), .IN2(n53), .QN(\ab[11][1] ) );
  NOR2X0 U312 ( .IN1(n33), .IN2(n53), .QN(\ab[11][15] ) );
  NOR2X0 U313 ( .IN1(n34), .IN2(n53), .QN(\ab[11][14] ) );
  NOR2X0 U314 ( .IN1(n35), .IN2(n53), .QN(\ab[11][13] ) );
  NOR2X0 U315 ( .IN1(n36), .IN2(n53), .QN(\ab[11][12] ) );
  NOR2X0 U316 ( .IN1(n37), .IN2(n53), .QN(\ab[11][11] ) );
  NOR2X0 U317 ( .IN1(n38), .IN2(n53), .QN(\ab[11][10] ) );
  NOR2X0 U318 ( .IN1(n48), .IN2(n53), .QN(\ab[11][0] ) );
  NOR2X0 U319 ( .IN1(n39), .IN2(n54), .QN(\ab[10][9] ) );
  NOR2X0 U320 ( .IN1(n40), .IN2(n54), .QN(\ab[10][8] ) );
  NOR2X0 U321 ( .IN1(n41), .IN2(n54), .QN(\ab[10][7] ) );
  NOR2X0 U322 ( .IN1(n42), .IN2(n54), .QN(\ab[10][6] ) );
  NOR2X0 U323 ( .IN1(n43), .IN2(n54), .QN(\ab[10][5] ) );
  NOR2X0 U324 ( .IN1(n44), .IN2(n54), .QN(\ab[10][4] ) );
  NOR2X0 U325 ( .IN1(n45), .IN2(n54), .QN(\ab[10][3] ) );
  NOR2X0 U326 ( .IN1(n46), .IN2(n54), .QN(\ab[10][2] ) );
  NOR2X0 U327 ( .IN1(n47), .IN2(n54), .QN(\ab[10][1] ) );
  NOR2X0 U328 ( .IN1(n33), .IN2(n54), .QN(\ab[10][15] ) );
  NOR2X0 U329 ( .IN1(n34), .IN2(n54), .QN(\ab[10][14] ) );
  NOR2X0 U330 ( .IN1(n35), .IN2(n54), .QN(\ab[10][13] ) );
  NOR2X0 U331 ( .IN1(n36), .IN2(n54), .QN(\ab[10][12] ) );
  NOR2X0 U332 ( .IN1(n37), .IN2(n54), .QN(\ab[10][11] ) );
  NOR2X0 U333 ( .IN1(n38), .IN2(n54), .QN(\ab[10][10] ) );
  NOR2X0 U334 ( .IN1(n48), .IN2(n54), .QN(\ab[10][0] ) );
  NOR2X0 U335 ( .IN1(n39), .IN2(n64), .QN(\ab[0][9] ) );
  NOR2X0 U336 ( .IN1(n40), .IN2(n64), .QN(\ab[0][8] ) );
  NOR2X0 U337 ( .IN1(n41), .IN2(n64), .QN(\ab[0][7] ) );
  NOR2X0 U338 ( .IN1(n42), .IN2(n64), .QN(\ab[0][6] ) );
  NOR2X0 U339 ( .IN1(n43), .IN2(n64), .QN(\ab[0][5] ) );
  NOR2X0 U340 ( .IN1(n44), .IN2(n64), .QN(\ab[0][4] ) );
  NOR2X0 U341 ( .IN1(n45), .IN2(n64), .QN(\ab[0][3] ) );
  NOR2X0 U342 ( .IN1(n46), .IN2(n64), .QN(\ab[0][2] ) );
  NOR2X0 U343 ( .IN1(n47), .IN2(n64), .QN(\ab[0][1] ) );
  NOR2X0 U344 ( .IN1(n33), .IN2(n64), .QN(\ab[0][15] ) );
  NOR2X0 U345 ( .IN1(n34), .IN2(n64), .QN(\ab[0][14] ) );
  NOR2X0 U346 ( .IN1(n35), .IN2(n64), .QN(\ab[0][13] ) );
  NOR2X0 U347 ( .IN1(n36), .IN2(n64), .QN(\ab[0][12] ) );
  NOR2X0 U348 ( .IN1(n37), .IN2(n64), .QN(\ab[0][11] ) );
  NOR2X0 U349 ( .IN1(n38), .IN2(n64), .QN(\ab[0][10] ) );
  NOR2X0 U350 ( .IN1(n48), .IN2(n64), .QN(PRODUCT[0]) );
endmodule


module betterNeighborsInMyCluster ( clock, nrst, en, start, address, wr_en, 
        data_in, MY_CLUSTER_ID, mybest, besthop, bestvalue, bestneighborID, 
        nextsinks, data_out, done );
  output [10:0] address;
  input [15:0] data_in;
  input [15:0] MY_CLUSTER_ID;
  input [15:0] mybest;
  output [15:0] besthop;
  output [15:0] bestvalue;
  output [15:0] bestneighborID;
  output [15:0] nextsinks;
  output [15:0] data_out;
  input clock, nrst, en, start;
  output wr_en, done;
  wire   N130, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N150, N151, N153, N154, N155, N156, N157,
         N158, N159, N160, N163, N164, N165, N166, N167, N168, N169, N170,
         N171, N172, N188, N189, N190, N191, N192, N193, N194, N230, N231,
         N232, N233, N234, N235, N236, N237, N267, N268, N269, N270, N271,
         N272, N273, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N330, N331, N332, N333, N334,
         N335, N336, N337, N338, N339, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N374, N375, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N406, N413, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N446, N447, N448, N449, N450, N451, N452,
         N453, N454, N455, N456, N457, N458, N459, N472, N473, N474, N475,
         N476, N477, N478, N479, N480, N481, N483, N486, N487, N488, N489,
         N490, N491, N492, N493, N494, N495, N496, N497, N498, N499, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N534,
         N535, N536, N537, N538, N539, N540, N1262, N1264, N1266, N1268, N1270,
         N1272, N1276, n55, n56, n57, n58, n59, n60, n61, n62, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, N317, N316, N315, N314, N313,
         N312, N311, N310, \add_218/carry[10] , \add_218/carry[9] ,
         \add_218/carry[8] , \add_218/carry[7] , \add_218/carry[6] ,
         \add_218/carry[5] , \add_212/carry[10] , \add_212/carry[9] ,
         \add_212/carry[8] , \add_212/carry[7] , \add_212/carry[6] ,
         \add_212/carry[5] , \add_199/carry[10] , \add_199/carry[9] ,
         \add_199/carry[8] , \add_199/carry[7] , \add_199/carry[6] ,
         \add_199/carry[5] , \add_177/carry[10] , \add_177/carry[9] ,
         \add_177/carry[8] , \add_177/carry[7] , \add_177/carry[6] ,
         \add_177/carry[5] , \add_137/carry[10] , \add_137/carry[9] ,
         \add_137/carry[8] , \add_137/carry[7] , \add_137/carry[6] ,
         \add_137/carry[5] , \add_128/carry[10] , \add_128/carry[9] ,
         \add_128/carry[8] , \add_128/carry[7] , \add_128/carry[6] ,
         \add_128/carry[5] , \add_117/carry[10] , \add_117/carry[9] ,
         \add_117/carry[8] , \add_117/carry[7] , \add_117/carry[6] ,
         \add_117/carry[5] , \add_108/carry[10] , \add_108/carry[9] ,
         \add_108/carry[8] , \add_108/carry[7] , \add_108/carry[6] ,
         \add_108/carry[5] , \r221/carry[10] , \r221/carry[9] ,
         \r221/carry[8] , \r221/carry[7] , \r221/carry[6] , \r221/carry[5] ,
         \r212/carry[10] , \r212/carry[9] , \r212/carry[8] , \r212/carry[7] ,
         \r212/carry[6] , \r212/carry[5] , \add_151/carry[10] ,
         \add_151/carry[9] , \add_151/carry[8] , \add_151/carry[7] ,
         \add_151/carry[6] , \add_151/carry[5] , n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990;
  wire   [3:0] state;
  wire   [15:0] i;
  wire   [15:0] neighborCount;
  wire   [15:0] betterneighborCount;
  wire   [30:0] fpTemp;
  wire   [15:0] j;
  wire   [15:0] k;
  wire   [15:0] batteryStat;
  wire   [15:0] knownSinkCount;
  wire   [15:0] neighborID;
  wire   [15:0] qValue;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;
  assign besthop[0] = N163;
  assign besthop[1] = N164;

  DFFX1 \fpTemp_reg[14]  ( .D(n395), .CLK(clock), .Q(n768), .QN(n984) );
  DFFX1 \fpTemp_reg[13]  ( .D(n394), .CLK(clock), .Q(n769), .QN(n983) );
  DFFX1 \fpTemp_reg[12]  ( .D(n393), .CLK(clock), .Q(n770), .QN(n982) );
  DFFX1 \fpTemp_reg[11]  ( .D(n392), .CLK(clock), .Q(n771), .QN(n981) );
  DFFX1 \fpTemp_reg[10]  ( .D(n391), .CLK(clock), .Q(n772), .QN(n980) );
  DFFX1 \fpTemp_reg[9]  ( .D(n390), .CLK(clock), .Q(n773), .QN(n979) );
  DFFX1 \fpTemp_reg[8]  ( .D(n389), .CLK(clock), .Q(n774), .QN(n978) );
  DFFX1 \fpTemp_reg[7]  ( .D(n388), .CLK(clock), .Q(n775), .QN(n977) );
  DFFX1 \fpTemp_reg[6]  ( .D(n387), .CLK(clock), .Q(n776), .QN(n976) );
  DFFX1 \fpTemp_reg[5]  ( .D(n386), .CLK(clock), .Q(n777), .QN(n975) );
  DFFX1 \fpTemp_reg[4]  ( .D(n385), .CLK(clock), .Q(n778), .QN(n974) );
  DFFX1 \fpTemp_reg[3]  ( .D(n384), .CLK(clock), .Q(n779), .QN(n973) );
  DFFX1 \fpTemp_reg[2]  ( .D(n383), .CLK(clock), .Q(n780), .QN(n972) );
  DFFX1 \fpTemp_reg[1]  ( .D(n382), .CLK(clock), .Q(n781), .QN(n971) );
  DFFX1 \fpTemp_reg[0]  ( .D(n381), .CLK(clock), .Q(n782), .QN(n989) );
  DFFX1 \bestvalue_buf_reg[9]  ( .D(n262), .CLK(clock), .Q(bestvalue[9]), .QN(
        n960) );
  DFFX1 \bestvalue_buf_reg[8]  ( .D(n263), .CLK(clock), .Q(bestvalue[8]), .QN(
        n961) );
  DFFX1 \bestvalue_buf_reg[7]  ( .D(n264), .CLK(clock), .Q(bestvalue[7]), .QN(
        n962) );
  DFFX1 \bestvalue_buf_reg[6]  ( .D(n265), .CLK(clock), .Q(bestvalue[6]), .QN(
        n963) );
  DFFX1 \bestvalue_buf_reg[5]  ( .D(n266), .CLK(clock), .Q(bestvalue[5]), .QN(
        n964) );
  DFFX1 \bestvalue_buf_reg[4]  ( .D(n267), .CLK(clock), .Q(bestvalue[4]), .QN(
        n965) );
  DFFX1 \bestvalue_buf_reg[3]  ( .D(n268), .CLK(clock), .Q(bestvalue[3]), .QN(
        n966) );
  DFFX1 \bestvalue_buf_reg[2]  ( .D(n269), .CLK(clock), .Q(bestvalue[2]), .QN(
        n967) );
  DFFX1 \bestvalue_buf_reg[1]  ( .D(n270), .CLK(clock), .Q(bestvalue[1]), .QN(
        n968) );
  DFFX1 \besthop_buf_reg[6]  ( .D(n291), .CLK(clock), .Q(besthop[6]), .QN(n969) );
  DFFX1 \besthop_buf_reg[0]  ( .D(n297), .CLK(clock), .Q(N163), .QN(n970) );
  betterNeighborsInMyCluster_DW01_inc_0 add_168 ( .A(fpTemp[30:15]), .SUM({
        N389, N388, N387, N386, N385, N384, N383, N382, N381, N380, N379, N378, 
        N377, N376, N375, N374}) );
  betterNeighborsInMyCluster_DW01_inc_1 add_146 ( .A(betterneighborCount), 
        .SUM({N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292}) );
  betterNeighborsInMyCluster_DW01_inc_2 r209 ( .A({i[15:2], N331, N330}), 
        .SUM({N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, N138, 
        N137, N136, N135, N151, N150}) );
  betterNeighborsInMyCluster_DW01_inc_3 add_211 ( .A({j[15:2], N473, N472}), 
        .SUM({N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N502, N501}) );
  betterNeighborsInMyCluster_DW02_mult_1 mult_163 ( .A({1'b1, 1'b0, 1'b1, 1'b0}), .B(batteryStat), .TC(1'b0), .PRODUCT({N371, N370, N369, N368, N367, N366, 
        N365, N364, N363, N362, N361, N360, N359, N358, N357, N356, N355, N354, 
        N353, SYNOPSYS_UNCONNECTED__0}) );
  betterNeighborsInMyCluster_DW02_mult_0 mult_184 ( .A(qValue), .B(data_in), 
        .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__1, N458, N457, N456, N455, 
        N454, N453, N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, 
        N442, N441, N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, 
        N430, N429, N428}) );
  DFFX1 done_buf_reg ( .D(n332), .CLK(clock), .Q(done) );
  DFFX1 \neighborCount_reg[15]  ( .D(n476), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n477), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n478), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n479), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n480), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n481), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n482), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n483), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n484), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n485), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n486), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n487), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n488), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n489), .CLK(clock), .Q(neighborCount[2])
         );
  DFFX1 \neighborCount_reg[1]  ( .D(n490), .CLK(clock), .Q(neighborCount[1]), 
        .QN(n622) );
  DFFX1 \neighborCount_reg[0]  ( .D(n527), .CLK(clock), .Q(neighborCount[0]), 
        .QN(n624) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n460), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n461), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n462), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n463), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n464), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n465), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n466), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n467), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n468), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n469), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n470), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n471), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n472), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n473), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n474), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n599) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n475), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n598) );
  DFFX1 \j_reg[15]  ( .D(n444), .CLK(clock), .Q(j[15]) );
  DFFX1 \j_reg[14]  ( .D(n445), .CLK(clock), .Q(j[14]) );
  DFFX1 \j_reg[13]  ( .D(n446), .CLK(clock), .Q(j[13]) );
  DFFX1 \j_reg[12]  ( .D(n447), .CLK(clock), .Q(j[12]) );
  DFFX1 \j_reg[11]  ( .D(n448), .CLK(clock), .Q(j[11]) );
  DFFX1 \j_reg[10]  ( .D(n449), .CLK(clock), .Q(j[10]) );
  DFFX1 \j_reg[9]  ( .D(n450), .CLK(clock), .Q(j[9]) );
  DFFX1 \j_reg[8]  ( .D(n451), .CLK(clock), .Q(j[8]) );
  DFFX1 \j_reg[7]  ( .D(n452), .CLK(clock), .Q(j[7]) );
  DFFX1 \j_reg[6]  ( .D(n453), .CLK(clock), .Q(j[6]) );
  DFFX1 \j_reg[5]  ( .D(n454), .CLK(clock), .Q(j[5]) );
  DFFX1 \j_reg[4]  ( .D(n455), .CLK(clock), .Q(j[4]) );
  DFFX1 \j_reg[3]  ( .D(n456), .CLK(clock), .Q(j[3]) );
  DFFX1 \j_reg[2]  ( .D(n457), .CLK(clock), .Q(j[2]), .QN(N474) );
  DFFX1 \j_reg[1]  ( .D(n458), .CLK(clock), .Q(N473) );
  DFFX1 \j_reg[0]  ( .D(n459), .CLK(clock), .Q(N472) );
  DFFX1 \batteryStat_reg[15]  ( .D(n507), .CLK(clock), .Q(batteryStat[15]) );
  DFFX1 \batteryStat_reg[14]  ( .D(n508), .CLK(clock), .Q(batteryStat[14]) );
  DFFX1 \batteryStat_reg[13]  ( .D(n509), .CLK(clock), .Q(batteryStat[13]) );
  DFFX1 \batteryStat_reg[12]  ( .D(n510), .CLK(clock), .Q(batteryStat[12]) );
  DFFX1 \batteryStat_reg[11]  ( .D(n511), .CLK(clock), .Q(batteryStat[11]) );
  DFFX1 \batteryStat_reg[10]  ( .D(n512), .CLK(clock), .Q(batteryStat[10]) );
  DFFX1 \batteryStat_reg[9]  ( .D(n513), .CLK(clock), .Q(batteryStat[9]) );
  DFFX1 \batteryStat_reg[8]  ( .D(n514), .CLK(clock), .Q(batteryStat[8]) );
  DFFX1 \batteryStat_reg[7]  ( .D(n515), .CLK(clock), .Q(batteryStat[7]) );
  DFFX1 \batteryStat_reg[6]  ( .D(n516), .CLK(clock), .Q(batteryStat[6]) );
  DFFX1 \batteryStat_reg[5]  ( .D(n517), .CLK(clock), .Q(batteryStat[5]) );
  DFFX1 \batteryStat_reg[4]  ( .D(n518), .CLK(clock), .Q(batteryStat[4]) );
  DFFX1 \batteryStat_reg[3]  ( .D(n519), .CLK(clock), .Q(batteryStat[3]) );
  DFFX1 \batteryStat_reg[2]  ( .D(n520), .CLK(clock), .Q(batteryStat[2]) );
  DFFX1 \batteryStat_reg[1]  ( .D(n521), .CLK(clock), .Q(batteryStat[1]) );
  DFFX1 \batteryStat_reg[0]  ( .D(n522), .CLK(clock), .Q(batteryStat[0]) );
  DFFX1 \neighborID_reg[15]  ( .D(n491), .CLK(clock), .Q(neighborID[15]) );
  DFFX1 \neighborID_reg[14]  ( .D(n492), .CLK(clock), .Q(neighborID[14]) );
  DFFX1 \neighborID_reg[13]  ( .D(n493), .CLK(clock), .Q(neighborID[13]) );
  DFFX1 \neighborID_reg[12]  ( .D(n494), .CLK(clock), .Q(neighborID[12]) );
  DFFX1 \neighborID_reg[11]  ( .D(n495), .CLK(clock), .Q(neighborID[11]) );
  DFFX1 \neighborID_reg[10]  ( .D(n496), .CLK(clock), .Q(neighborID[10]) );
  DFFX1 \neighborID_reg[9]  ( .D(n497), .CLK(clock), .Q(neighborID[9]) );
  DFFX1 \neighborID_reg[8]  ( .D(n498), .CLK(clock), .Q(neighborID[8]) );
  DFFX1 \neighborID_reg[7]  ( .D(n499), .CLK(clock), .Q(neighborID[7]) );
  DFFX1 \neighborID_reg[6]  ( .D(n500), .CLK(clock), .Q(neighborID[6]) );
  DFFX1 \neighborID_reg[5]  ( .D(n501), .CLK(clock), .Q(neighborID[5]) );
  DFFX1 \neighborID_reg[4]  ( .D(n502), .CLK(clock), .Q(neighborID[4]) );
  DFFX1 \neighborID_reg[3]  ( .D(n503), .CLK(clock), .Q(neighborID[3]) );
  DFFX1 \neighborID_reg[2]  ( .D(n504), .CLK(clock), .Q(neighborID[2]) );
  DFFX1 \neighborID_reg[1]  ( .D(n505), .CLK(clock), .Q(neighborID[1]), .QN(
        n686) );
  DFFX1 \neighborID_reg[0]  ( .D(n506), .CLK(clock), .Q(neighborID[0]) );
  DFFX1 \bestneighborID_buf_reg[15]  ( .D(n364), .CLK(clock), .Q(
        bestneighborID[15]) );
  DFFX1 \bestneighborID_buf_reg[14]  ( .D(n363), .CLK(clock), .Q(
        bestneighborID[14]) );
  DFFX1 \bestneighborID_buf_reg[13]  ( .D(n362), .CLK(clock), .Q(
        bestneighborID[13]) );
  DFFX1 \bestneighborID_buf_reg[12]  ( .D(n361), .CLK(clock), .Q(
        bestneighborID[12]) );
  DFFX1 \bestneighborID_buf_reg[0]  ( .D(n349), .CLK(clock), .Q(
        bestneighborID[0]) );
  DFFX1 \k_reg[15]  ( .D(n380), .CLK(clock), .Q(k[15]) );
  DFFX1 \k_reg[14]  ( .D(n365), .CLK(clock), .Q(k[14]) );
  DFFX1 \k_reg[13]  ( .D(n366), .CLK(clock), .Q(k[13]) );
  DFFX1 \k_reg[12]  ( .D(n367), .CLK(clock), .Q(k[12]) );
  DFFX1 \k_reg[11]  ( .D(n368), .CLK(clock), .Q(k[11]) );
  DFFX1 \k_reg[10]  ( .D(n369), .CLK(clock), .Q(k[10]) );
  DFFX1 \state_reg[0]  ( .D(n525), .CLK(clock), .Q(state[0]), .QN(n952) );
  DFFX1 \state_reg[1]  ( .D(n524), .CLK(clock), .Q(state[1]), .QN(n897) );
  DFFX1 \nextsinks_buf_reg[6]  ( .D(n421), .CLK(clock), .Q(nextsinks[6]) );
  DFFX1 \nextsinks_buf_reg[0]  ( .D(n427), .CLK(clock), .Q(nextsinks[0]) );
  DFFX1 \bestneighborID_buf_reg[11]  ( .D(n360), .CLK(clock), .Q(
        bestneighborID[11]) );
  DFFX1 \bestneighborID_buf_reg[10]  ( .D(n359), .CLK(clock), .Q(
        bestneighborID[10]) );
  DFFX1 \bestneighborID_buf_reg[9]  ( .D(n358), .CLK(clock), .Q(
        bestneighborID[9]) );
  DFFX1 \bestneighborID_buf_reg[8]  ( .D(n357), .CLK(clock), .Q(
        bestneighborID[8]) );
  DFFX1 \bestneighborID_buf_reg[7]  ( .D(n356), .CLK(clock), .Q(
        bestneighborID[7]) );
  DFFX1 \bestneighborID_buf_reg[6]  ( .D(n355), .CLK(clock), .Q(
        bestneighborID[6]) );
  DFFX1 \bestneighborID_buf_reg[5]  ( .D(n354), .CLK(clock), .Q(
        bestneighborID[5]) );
  DFFX1 \bestneighborID_buf_reg[4]  ( .D(n353), .CLK(clock), .Q(
        bestneighborID[4]) );
  DFFX1 \bestneighborID_buf_reg[3]  ( .D(n352), .CLK(clock), .Q(
        bestneighborID[3]) );
  DFFX1 \bestneighborID_buf_reg[2]  ( .D(n351), .CLK(clock), .Q(
        bestneighborID[2]) );
  DFFX1 \bestneighborID_buf_reg[1]  ( .D(n350), .CLK(clock), .Q(
        bestneighborID[1]) );
  DFFX1 \nextsinks_buf_reg[15]  ( .D(n412), .CLK(clock), .Q(nextsinks[15]) );
  DFFX1 \nextsinks_buf_reg[14]  ( .D(n413), .CLK(clock), .Q(nextsinks[14]) );
  DFFX1 \nextsinks_buf_reg[13]  ( .D(n414), .CLK(clock), .Q(nextsinks[13]) );
  DFFX1 \nextsinks_buf_reg[12]  ( .D(n415), .CLK(clock), .Q(nextsinks[12]) );
  DFFX1 \nextsinks_buf_reg[11]  ( .D(n416), .CLK(clock), .Q(nextsinks[11]) );
  DFFX1 \nextsinks_buf_reg[10]  ( .D(n417), .CLK(clock), .Q(nextsinks[10]) );
  DFFX1 \nextsinks_buf_reg[9]  ( .D(n418), .CLK(clock), .Q(nextsinks[9]) );
  DFFX1 \nextsinks_buf_reg[8]  ( .D(n419), .CLK(clock), .Q(nextsinks[8]) );
  DFFX1 \nextsinks_buf_reg[7]  ( .D(n420), .CLK(clock), .Q(nextsinks[7]) );
  DFFX1 \nextsinks_buf_reg[5]  ( .D(n422), .CLK(clock), .Q(nextsinks[5]) );
  DFFX1 \nextsinks_buf_reg[4]  ( .D(n423), .CLK(clock), .Q(nextsinks[4]) );
  DFFX1 \nextsinks_buf_reg[3]  ( .D(n424), .CLK(clock), .Q(nextsinks[3]) );
  DFFX1 \nextsinks_buf_reg[2]  ( .D(n425), .CLK(clock), .Q(nextsinks[2]) );
  DFFX1 \nextsinks_buf_reg[1]  ( .D(n426), .CLK(clock), .Q(nextsinks[1]) );
  DFFX1 \state_reg[2]  ( .D(n523), .CLK(clock), .Q(state[2]), .QN(n935) );
  DFFX1 \state_reg[3]  ( .D(n526), .CLK(clock), .Q(state[3]), .QN(n951) );
  DFFX1 \address_count_reg[8]  ( .D(n279), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[5]  ( .D(n282), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n283), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[10]  ( .D(n277), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n278), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[7]  ( .D(n280), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[3]  ( .D(n284), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[6]  ( .D(n281), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[2]  ( .D(n285), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[1]  ( .D(n286), .CLK(clock), .Q(address[1]) );
  DFFX1 wr_en_buf_reg ( .D(n331), .CLK(clock), .Q(wr_en) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n299), .CLK(clock), .Q(data_out[15]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n300), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n301), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n302), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n303), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n304), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n305), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n306), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n307), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n308), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n309), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n310), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n311), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n312), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n313), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n314), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \qValue_reg[0]  ( .D(n333), .CLK(clock), .Q(qValue[0]) );
  DFFX1 \qValue_reg[1]  ( .D(n334), .CLK(clock), .Q(qValue[1]) );
  DFFX1 \qValue_reg[2]  ( .D(n335), .CLK(clock), .Q(qValue[2]) );
  DFFX1 \qValue_reg[3]  ( .D(n336), .CLK(clock), .Q(qValue[3]) );
  DFFX1 \qValue_reg[4]  ( .D(n337), .CLK(clock), .Q(qValue[4]) );
  DFFX1 \qValue_reg[5]  ( .D(n338), .CLK(clock), .Q(qValue[5]) );
  DFFX1 \qValue_reg[6]  ( .D(n339), .CLK(clock), .Q(qValue[6]) );
  DFFX1 \qValue_reg[7]  ( .D(n340), .CLK(clock), .Q(qValue[7]) );
  DFFX1 \qValue_reg[8]  ( .D(n341), .CLK(clock), .Q(qValue[8]) );
  DFFX1 \qValue_reg[9]  ( .D(n342), .CLK(clock), .Q(qValue[9]) );
  DFFX1 \qValue_reg[10]  ( .D(n343), .CLK(clock), .Q(qValue[10]) );
  DFFX1 \qValue_reg[11]  ( .D(n344), .CLK(clock), .Q(qValue[11]) );
  DFFX1 \qValue_reg[12]  ( .D(n345), .CLK(clock), .Q(qValue[12]) );
  DFFX1 \qValue_reg[13]  ( .D(n346), .CLK(clock), .Q(qValue[13]) );
  DFFX1 \qValue_reg[14]  ( .D(n347), .CLK(clock), .Q(qValue[14]) );
  DFFX1 \qValue_reg[15]  ( .D(n348), .CLK(clock), .Q(qValue[15]) );
  DFFX1 \bestvalue_buf_reg[0]  ( .D(n298), .CLK(clock), .Q(bestvalue[0]), .QN(
        n648) );
  DFFX1 \besthop_buf_reg[15]  ( .D(n271), .CLK(clock), .Q(besthop[15]) );
  DFFX1 \besthop_buf_reg[14]  ( .D(n272), .CLK(clock), .Q(besthop[14]) );
  DFFX1 \besthop_buf_reg[13]  ( .D(n273), .CLK(clock), .Q(besthop[13]) );
  DFFX1 \besthop_buf_reg[12]  ( .D(n274), .CLK(clock), .Q(besthop[12]) );
  DFFX1 \besthop_buf_reg[11]  ( .D(n275), .CLK(clock), .Q(besthop[11]) );
  DFFX1 \besthop_buf_reg[10]  ( .D(n276), .CLK(clock), .Q(besthop[10]) );
  DFFX1 \besthop_buf_reg[9]  ( .D(n288), .CLK(clock), .Q(besthop[9]) );
  DFFX1 \besthop_buf_reg[8]  ( .D(n289), .CLK(clock), .Q(besthop[8]) );
  DFFX1 \besthop_buf_reg[7]  ( .D(n290), .CLK(clock), .Q(besthop[7]) );
  DFFX1 \besthop_buf_reg[5]  ( .D(n292), .CLK(clock), .Q(besthop[5]) );
  DFFX1 \besthop_buf_reg[4]  ( .D(n293), .CLK(clock), .Q(besthop[4]) );
  DFFX1 \besthop_buf_reg[3]  ( .D(n294), .CLK(clock), .Q(besthop[3]) );
  DFFX1 \besthop_buf_reg[2]  ( .D(n295), .CLK(clock), .Q(besthop[2]), .QN(N165) );
  DFFX1 \besthop_buf_reg[1]  ( .D(n296), .CLK(clock), .Q(N164) );
  DFFX1 \k_reg[9]  ( .D(n370), .CLK(clock), .Q(k[9]), .QN(n55) );
  DFFX1 \k_reg[8]  ( .D(n371), .CLK(clock), .Q(k[8]), .QN(n56) );
  DFFX1 \k_reg[7]  ( .D(n372), .CLK(clock), .Q(k[7]), .QN(n57) );
  DFFX1 \k_reg[6]  ( .D(n373), .CLK(clock), .Q(k[6]), .QN(n58) );
  DFFX1 \k_reg[5]  ( .D(n374), .CLK(clock), .Q(k[5]), .QN(n59) );
  DFFX1 \k_reg[4]  ( .D(n375), .CLK(clock), .Q(k[4]), .QN(n60) );
  DFFX1 \k_reg[2]  ( .D(n377), .CLK(clock), .Q(k[2]), .QN(n61) );
  DFFX1 \k_reg[0]  ( .D(n379), .CLK(clock), .Q(k[0]), .QN(n62) );
  DFFX1 \k_reg[3]  ( .D(n376), .CLK(clock), .Q(k[3]), .QN(n988) );
  DFFX1 \k_reg[1]  ( .D(n378), .CLK(clock), .Q(k[1]), .QN(n987) );
  DFFX1 \address_count_reg[0]  ( .D(n287), .CLK(clock), .Q(address[0]), .QN(
        n990) );
  DFFX1 \i_reg[15]  ( .D(n443), .CLK(clock), .Q(i[15]) );
  DFFX1 \i_reg[14]  ( .D(n428), .CLK(clock), .Q(i[14]) );
  DFFX1 \i_reg[13]  ( .D(n429), .CLK(clock), .Q(i[13]) );
  DFFX1 \i_reg[12]  ( .D(n430), .CLK(clock), .Q(i[12]) );
  DFFX1 \i_reg[11]  ( .D(n431), .CLK(clock), .Q(i[11]) );
  DFFX1 \i_reg[10]  ( .D(n432), .CLK(clock), .Q(i[10]) );
  DFFX1 \i_reg[9]  ( .D(n433), .CLK(clock), .Q(i[9]) );
  DFFX1 \i_reg[8]  ( .D(n434), .CLK(clock), .Q(i[8]) );
  DFFX1 \i_reg[7]  ( .D(n435), .CLK(clock), .Q(i[7]) );
  DFFX1 \i_reg[6]  ( .D(n436), .CLK(clock), .Q(i[6]), .QN(n985) );
  DFFX1 \i_reg[5]  ( .D(n437), .CLK(clock), .Q(i[5]) );
  DFFX1 \i_reg[4]  ( .D(n438), .CLK(clock), .Q(i[4]) );
  DFFX1 \i_reg[3]  ( .D(n439), .CLK(clock), .Q(i[3]) );
  DFFX1 \i_reg[2]  ( .D(n440), .CLK(clock), .Q(i[2]), .QN(N332) );
  DFFX1 \i_reg[1]  ( .D(n441), .CLK(clock), .Q(N331) );
  DFFX1 \i_reg[0]  ( .D(n442), .CLK(clock), .Q(N330), .QN(n986) );
  DFFX1 \betterneighborCount_reg[15]  ( .D(n315), .CLK(clock), .Q(
        betterneighborCount[15]) );
  DFFX1 \betterneighborCount_reg[14]  ( .D(n316), .CLK(clock), .Q(
        betterneighborCount[14]) );
  DFFX1 \betterneighborCount_reg[13]  ( .D(n317), .CLK(clock), .Q(
        betterneighborCount[13]) );
  DFFX1 \betterneighborCount_reg[12]  ( .D(n318), .CLK(clock), .Q(
        betterneighborCount[12]) );
  DFFX1 \betterneighborCount_reg[11]  ( .D(n319), .CLK(clock), .Q(
        betterneighborCount[11]) );
  DFFX1 \betterneighborCount_reg[10]  ( .D(n320), .CLK(clock), .Q(
        betterneighborCount[10]) );
  DFFX1 \betterneighborCount_reg[9]  ( .D(n321), .CLK(clock), .Q(
        betterneighborCount[9]) );
  DFFX1 \betterneighborCount_reg[8]  ( .D(n322), .CLK(clock), .Q(
        betterneighborCount[8]) );
  DFFX1 \betterneighborCount_reg[7]  ( .D(n323), .CLK(clock), .Q(
        betterneighborCount[7]) );
  DFFX1 \betterneighborCount_reg[6]  ( .D(n324), .CLK(clock), .Q(
        betterneighborCount[6]) );
  DFFX1 \betterneighborCount_reg[5]  ( .D(n325), .CLK(clock), .Q(
        betterneighborCount[5]) );
  DFFX1 \betterneighborCount_reg[4]  ( .D(n326), .CLK(clock), .Q(
        betterneighborCount[4]) );
  DFFX1 \betterneighborCount_reg[3]  ( .D(n327), .CLK(clock), .Q(
        betterneighborCount[3]) );
  DFFX1 \betterneighborCount_reg[2]  ( .D(n328), .CLK(clock), .Q(
        betterneighborCount[2]) );
  DFFX1 \betterneighborCount_reg[1]  ( .D(n329), .CLK(clock), .Q(
        betterneighborCount[1]) );
  DFFX1 \betterneighborCount_reg[0]  ( .D(n330), .CLK(clock), .Q(
        betterneighborCount[0]) );
  DFFX1 \fpTemp_reg[15]  ( .D(n396), .CLK(clock), .Q(fpTemp[15]) );
  DFFX1 \fpTemp_reg[16]  ( .D(n397), .CLK(clock), .Q(fpTemp[16]) );
  DFFX1 \fpTemp_reg[17]  ( .D(n398), .CLK(clock), .Q(fpTemp[17]) );
  DFFX1 \fpTemp_reg[18]  ( .D(n399), .CLK(clock), .Q(fpTemp[18]) );
  DFFX1 \fpTemp_reg[19]  ( .D(n400), .CLK(clock), .Q(fpTemp[19]) );
  DFFX1 \fpTemp_reg[20]  ( .D(n401), .CLK(clock), .Q(fpTemp[20]) );
  DFFX1 \fpTemp_reg[21]  ( .D(n402), .CLK(clock), .Q(fpTemp[21]) );
  DFFX1 \fpTemp_reg[22]  ( .D(n403), .CLK(clock), .Q(fpTemp[22]) );
  DFFX1 \fpTemp_reg[23]  ( .D(n404), .CLK(clock), .Q(fpTemp[23]) );
  DFFX1 \fpTemp_reg[24]  ( .D(n405), .CLK(clock), .Q(fpTemp[24]) );
  DFFX1 \fpTemp_reg[25]  ( .D(n406), .CLK(clock), .Q(fpTemp[25]) );
  DFFX1 \fpTemp_reg[26]  ( .D(n407), .CLK(clock), .Q(fpTemp[26]) );
  DFFX1 \fpTemp_reg[27]  ( .D(n408), .CLK(clock), .Q(fpTemp[27]) );
  DFFX1 \fpTemp_reg[28]  ( .D(n409), .CLK(clock), .Q(fpTemp[28]) );
  DFFX1 \fpTemp_reg[29]  ( .D(n410), .CLK(clock), .Q(fpTemp[29]) );
  DFFX1 \fpTemp_reg[30]  ( .D(n411), .CLK(clock), .Q(fpTemp[30]) );
  DFFX1 \bestvalue_buf_reg[15]  ( .D(n256), .CLK(clock), .Q(bestvalue[15]), 
        .QN(n954) );
  DFFX1 \bestvalue_buf_reg[14]  ( .D(n257), .CLK(clock), .Q(bestvalue[14]), 
        .QN(n955) );
  DFFX1 \bestvalue_buf_reg[13]  ( .D(n258), .CLK(clock), .Q(bestvalue[13]), 
        .QN(n956) );
  DFFX1 \bestvalue_buf_reg[12]  ( .D(n259), .CLK(clock), .Q(bestvalue[12]), 
        .QN(n957) );
  DFFX1 \bestvalue_buf_reg[11]  ( .D(n260), .CLK(clock), .Q(bestvalue[11]), 
        .QN(n958) );
  DFFX1 \bestvalue_buf_reg[10]  ( .D(n261), .CLK(clock), .Q(bestvalue[10]), 
        .QN(n959) );
  OR2X1 U516 ( .IN1(n736), .IN2(n741), .Q(n528) );
  OR2X1 U517 ( .IN1(n783), .IN2(n734), .Q(n529) );
  INVX0 U518 ( .INP(N446), .ZN(n653) );
  INVX0 U519 ( .INP(N452), .ZN(n659) );
  INVX0 U520 ( .INP(N450), .ZN(n657) );
  INVX0 U521 ( .INP(N447), .ZN(n654) );
  INVX0 U522 ( .INP(N449), .ZN(n656) );
  INVX0 U523 ( .INP(N453), .ZN(n660) );
  INVX0 U524 ( .INP(N455), .ZN(n662) );
  INVX0 U525 ( .INP(n529), .ZN(n534) );
  INVX0 U526 ( .INP(n529), .ZN(n535) );
  INVX0 U527 ( .INP(N444), .ZN(n651) );
  NOR2X0 U528 ( .IN1(n783), .IN2(n818), .QN(n805) );
  INVX0 U529 ( .INP(n709), .ZN(n836) );
  INVX0 U530 ( .INP(N443), .ZN(n650) );
  INVX0 U531 ( .INP(n819), .ZN(n815) );
  INVX0 U532 ( .INP(n691), .ZN(n837) );
  NOR2X0 U533 ( .IN1(n698), .IN2(N160), .QN(n834) );
  NOR2X0 U534 ( .IN1(n725), .IN2(N130), .QN(n737) );
  INVX0 U535 ( .INP(n702), .ZN(n835) );
  NOR2X0 U536 ( .IN1(n804), .IN2(n801), .QN(n803) );
  INVX0 U537 ( .INP(n763), .ZN(n764) );
  INVX0 U538 ( .INP(n528), .ZN(n532) );
  INVX0 U539 ( .INP(n528), .ZN(n530) );
  INVX0 U540 ( .INP(n528), .ZN(n531) );
  INVX0 U541 ( .INP(n528), .ZN(n533) );
  NOR2X0 U542 ( .IN1(n727), .IN2(N160), .QN(n838) );
  NOR2X0 U543 ( .IN1(n714), .IN2(N511), .QN(n754) );
  INVX0 U544 ( .INP(n542), .ZN(n550) );
  INVX0 U545 ( .INP(n537), .ZN(n545) );
  INVX0 U546 ( .INP(n538), .ZN(n546) );
  INVX0 U547 ( .INP(n539), .ZN(n547) );
  INVX0 U548 ( .INP(n540), .ZN(n548) );
  INVX0 U549 ( .INP(n541), .ZN(n549) );
  INVX0 U550 ( .INP(n536), .ZN(n544) );
  INVX0 U551 ( .INP(n696), .ZN(n802) );
  INVX0 U552 ( .INP(n745), .ZN(n746) );
  INVX0 U553 ( .INP(n695), .ZN(n738) );
  NAND2X1 U554 ( .IN1(n824), .IN2(n762), .QN(n823) );
  AND2X1 U555 ( .IN1(n824), .IN2(n532), .Q(n821) );
  INVX0 U556 ( .INP(n824), .ZN(n820) );
  NOR2X0 U557 ( .IN1(n813), .IN2(n816), .QN(n817) );
  NOR2X0 U558 ( .IN1(n813), .IN2(n811), .QN(n814) );
  NOR2X0 U559 ( .IN1(n742), .IN2(n815), .QN(n811) );
  INVX0 U560 ( .INP(n718), .ZN(n816) );
  NOR2X0 U561 ( .IN1(n802), .IN2(n742), .QN(n801) );
  NOR2X0 U562 ( .IN1(n696), .IN2(n741), .QN(n800) );
  NOR2X0 U563 ( .IN1(n708), .IN2(n741), .QN(n750) );
  NOR2X0 U564 ( .IN1(n759), .IN2(n742), .QN(n756) );
  NOR2X0 U565 ( .IN1(n724), .IN2(n741), .QN(n740) );
  NOR2X0 U566 ( .IN1(n755), .IN2(n742), .QN(n752) );
  NOR2X0 U567 ( .IN1(n746), .IN2(n742), .QN(n743) );
  NOR2X0 U568 ( .IN1(n707), .IN2(n742), .QN(n739) );
  NOR2X0 U569 ( .IN1(n751), .IN2(n742), .QN(n749) );
  NOR2X0 U570 ( .IN1(n748), .IN2(n742), .QN(n687) );
  NOR2X0 U571 ( .IN1(n745), .IN2(n741), .QN(n744) );
  NOR2X0 U572 ( .IN1(n741), .IN2(n747), .QN(n688) );
  NOR2X0 U573 ( .IN1(n726), .IN2(n741), .QN(n767) );
  INVX0 U574 ( .INP(n813), .ZN(n806) );
  AND3X1 U575 ( .IN1(n697), .IN2(n791), .IN3(n792), .Q(n785) );
  NOR3X0 U576 ( .IN1(n741), .IN2(n790), .IN3(n697), .QN(n786) );
  NOR3X0 U577 ( .IN1(n756), .IN2(n758), .IN3(n741), .QN(n757) );
  NOR3X0 U578 ( .IN1(n697), .IN2(n741), .IN3(n793), .QN(n784) );
  INVX0 U579 ( .INP(N151), .ZN(n623) );
  INVX0 U580 ( .INP(N502), .ZN(n597) );
  INVX0 U581 ( .INP(N1276), .ZN(N420) );
  INVX0 U582 ( .INP(N486), .ZN(N503) );
  INVX0 U583 ( .INP(N442), .ZN(n649) );
  INVX0 U584 ( .INP(N451), .ZN(n658) );
  INVX0 U585 ( .INP(N445), .ZN(n652) );
  INVX0 U586 ( .INP(N448), .ZN(n655) );
  INVX0 U587 ( .INP(N454), .ZN(n661) );
  OA21X1 U588 ( .IN1(N459), .IN2(n742), .IN3(n783), .Q(n824) );
  INVX0 U589 ( .INP(N456), .ZN(n663) );
  INVX0 U590 ( .INP(N135), .ZN(N230) );
  INVX0 U591 ( .INP(N292), .ZN(N319) );
  INVX0 U592 ( .INP(N310), .ZN(N321) );
  AND2X1 U593 ( .IN1(n754), .IN2(nrst), .Q(n753) );
  AND2X1 U594 ( .IN1(n760), .IN2(nrst), .Q(n765) );
  INVX0 U595 ( .INP(MY_CLUSTER_ID[1]), .ZN(n574) );
  INVX0 U596 ( .INP(MY_CLUSTER_ID[0]), .ZN(n573) );
  INVX0 U597 ( .INP(nrst), .ZN(n741) );
  XOR2X1 U598 ( .IN1(i[9]), .IN2(\add_117/carry[10] ), .Q(N194) );
  XOR2X1 U599 ( .IN1(N493), .IN2(\add_212/carry[10] ), .Q(N510) );
  XOR2X1 U600 ( .IN1(besthop[9]), .IN2(\r212/carry[10] ), .Q(N172) );
  XNOR2X1 U601 ( .IN1(N317), .IN2(\add_151/carry[10] ), .Q(N328) );
  XOR2X1 U602 ( .IN1(N142), .IN2(\add_108/carry[10] ), .Q(N159) );
  XOR2X1 U603 ( .IN1(i[9]), .IN2(\add_137/carry[10] ), .Q(N273) );
  XNOR2X1 U604 ( .IN1(N1262), .IN2(\add_177/carry[10] ), .Q(N427) );
  XOR2X1 U605 ( .IN1(j[9]), .IN2(\add_199/carry[10] ), .Q(N481) );
  XOR2X1 U606 ( .IN1(N142), .IN2(\add_128/carry[10] ), .Q(N237) );
  XOR2X1 U607 ( .IN1(i[9]), .IN2(\r221/carry[10] ), .Q(N339) );
  XOR2X1 U608 ( .IN1(N142), .IN2(\add_218/carry[10] ), .Q(N540) );
  AND2X1 U609 ( .IN1(\add_117/carry[9] ), .IN2(i[8]), .Q(\add_117/carry[10] )
         );
  XOR2X1 U610 ( .IN1(i[8]), .IN2(\add_117/carry[9] ), .Q(N193) );
  AND2X1 U611 ( .IN1(\add_212/carry[9] ), .IN2(N492), .Q(\add_212/carry[10] )
         );
  XOR2X1 U612 ( .IN1(N492), .IN2(\add_212/carry[9] ), .Q(N509) );
  AND2X1 U613 ( .IN1(\r212/carry[9] ), .IN2(besthop[8]), .Q(\r212/carry[10] )
         );
  XOR2X1 U614 ( .IN1(besthop[8]), .IN2(\r212/carry[9] ), .Q(N171) );
  OR2X1 U615 ( .IN1(N316), .IN2(\add_151/carry[9] ), .Q(\add_151/carry[10] )
         );
  XNOR2X1 U616 ( .IN1(\add_151/carry[9] ), .IN2(N316), .Q(N327) );
  AND2X1 U617 ( .IN1(\add_108/carry[9] ), .IN2(N141), .Q(\add_108/carry[10] )
         );
  XOR2X1 U618 ( .IN1(N141), .IN2(\add_108/carry[9] ), .Q(N158) );
  AND2X1 U619 ( .IN1(\add_137/carry[9] ), .IN2(i[8]), .Q(\add_137/carry[10] )
         );
  XOR2X1 U620 ( .IN1(i[8]), .IN2(\add_137/carry[9] ), .Q(N272) );
  OR2X1 U621 ( .IN1(N1264), .IN2(\add_177/carry[9] ), .Q(\add_177/carry[10] )
         );
  XNOR2X1 U622 ( .IN1(\add_177/carry[9] ), .IN2(N1264), .Q(N426) );
  AND2X1 U623 ( .IN1(\add_199/carry[9] ), .IN2(j[8]), .Q(\add_199/carry[10] )
         );
  XOR2X1 U624 ( .IN1(j[8]), .IN2(\add_199/carry[9] ), .Q(N480) );
  AND2X1 U625 ( .IN1(\add_128/carry[9] ), .IN2(N141), .Q(\add_128/carry[10] )
         );
  XOR2X1 U626 ( .IN1(N141), .IN2(\add_128/carry[9] ), .Q(N236) );
  AND2X1 U627 ( .IN1(\r221/carry[9] ), .IN2(i[8]), .Q(\r221/carry[10] ) );
  XOR2X1 U628 ( .IN1(i[8]), .IN2(\r221/carry[9] ), .Q(N338) );
  AND2X1 U629 ( .IN1(\add_218/carry[9] ), .IN2(N141), .Q(\add_218/carry[10] )
         );
  XOR2X1 U630 ( .IN1(N141), .IN2(\add_218/carry[9] ), .Q(N539) );
  OR2X1 U631 ( .IN1(i[7]), .IN2(\add_117/carry[8] ), .Q(\add_117/carry[9] ) );
  XNOR2X1 U632 ( .IN1(\add_117/carry[8] ), .IN2(i[7]), .Q(N192) );
  AND2X1 U633 ( .IN1(\add_212/carry[8] ), .IN2(N491), .Q(\add_212/carry[9] )
         );
  XOR2X1 U634 ( .IN1(N491), .IN2(\add_212/carry[8] ), .Q(N508) );
  AND2X1 U635 ( .IN1(\r212/carry[8] ), .IN2(besthop[7]), .Q(\r212/carry[9] )
         );
  XOR2X1 U636 ( .IN1(besthop[7]), .IN2(\r212/carry[8] ), .Q(N170) );
  AND2X1 U637 ( .IN1(\add_151/carry[8] ), .IN2(N315), .Q(\add_151/carry[9] )
         );
  XOR2X1 U638 ( .IN1(N315), .IN2(\add_151/carry[8] ), .Q(N326) );
  AND2X1 U639 ( .IN1(\add_108/carry[8] ), .IN2(N140), .Q(\add_108/carry[9] )
         );
  XOR2X1 U640 ( .IN1(N140), .IN2(\add_108/carry[8] ), .Q(N157) );
  OR2X1 U641 ( .IN1(i[7]), .IN2(\add_137/carry[8] ), .Q(\add_137/carry[9] ) );
  XNOR2X1 U642 ( .IN1(\add_137/carry[8] ), .IN2(i[7]), .Q(N271) );
  AND2X1 U643 ( .IN1(\add_199/carry[8] ), .IN2(j[7]), .Q(\add_199/carry[9] )
         );
  XOR2X1 U644 ( .IN1(j[7]), .IN2(\add_199/carry[8] ), .Q(N479) );
  AND2X1 U645 ( .IN1(\add_177/carry[8] ), .IN2(N1266), .Q(\add_177/carry[9] )
         );
  XOR2X1 U646 ( .IN1(N1266), .IN2(\add_177/carry[8] ), .Q(N425) );
  AND2X1 U647 ( .IN1(\add_128/carry[8] ), .IN2(N140), .Q(\add_128/carry[9] )
         );
  XOR2X1 U648 ( .IN1(N140), .IN2(\add_128/carry[8] ), .Q(N235) );
  AND2X1 U649 ( .IN1(\r221/carry[8] ), .IN2(i[7]), .Q(\r221/carry[9] ) );
  XOR2X1 U650 ( .IN1(i[7]), .IN2(\r221/carry[8] ), .Q(N337) );
  AND2X1 U651 ( .IN1(\add_218/carry[8] ), .IN2(N140), .Q(\add_218/carry[9] )
         );
  XOR2X1 U652 ( .IN1(N140), .IN2(\add_218/carry[8] ), .Q(N538) );
  AND2X1 U653 ( .IN1(\add_117/carry[7] ), .IN2(i[6]), .Q(\add_117/carry[8] )
         );
  XOR2X1 U654 ( .IN1(i[6]), .IN2(\add_117/carry[7] ), .Q(N191) );
  AND2X1 U655 ( .IN1(\add_212/carry[7] ), .IN2(N490), .Q(\add_212/carry[8] )
         );
  XOR2X1 U656 ( .IN1(N490), .IN2(\add_212/carry[7] ), .Q(N507) );
  AND2X1 U657 ( .IN1(\r212/carry[7] ), .IN2(besthop[6]), .Q(\r212/carry[8] )
         );
  XOR2X1 U658 ( .IN1(besthop[6]), .IN2(\r212/carry[7] ), .Q(N169) );
  OR2X1 U659 ( .IN1(N139), .IN2(\add_108/carry[7] ), .Q(\add_108/carry[8] ) );
  XNOR2X1 U660 ( .IN1(\add_108/carry[7] ), .IN2(N139), .Q(N156) );
  AND2X1 U661 ( .IN1(\add_151/carry[7] ), .IN2(N314), .Q(\add_151/carry[8] )
         );
  XOR2X1 U662 ( .IN1(N314), .IN2(\add_151/carry[7] ), .Q(N325) );
  OR2X1 U663 ( .IN1(i[6]), .IN2(\add_137/carry[7] ), .Q(\add_137/carry[8] ) );
  XNOR2X1 U664 ( .IN1(\add_137/carry[7] ), .IN2(i[6]), .Q(N270) );
  AND2X1 U665 ( .IN1(\add_177/carry[7] ), .IN2(N1268), .Q(\add_177/carry[8] )
         );
  XOR2X1 U666 ( .IN1(N1268), .IN2(\add_177/carry[7] ), .Q(N424) );
  AND2X1 U667 ( .IN1(\add_199/carry[7] ), .IN2(j[6]), .Q(\add_199/carry[8] )
         );
  XOR2X1 U668 ( .IN1(j[6]), .IN2(\add_199/carry[7] ), .Q(N478) );
  OR2X1 U669 ( .IN1(N139), .IN2(\add_128/carry[7] ), .Q(\add_128/carry[8] ) );
  XNOR2X1 U670 ( .IN1(\add_128/carry[7] ), .IN2(N139), .Q(N234) );
  AND2X1 U671 ( .IN1(\r221/carry[7] ), .IN2(i[6]), .Q(\r221/carry[8] ) );
  XOR2X1 U672 ( .IN1(i[6]), .IN2(\r221/carry[7] ), .Q(N336) );
  OR2X1 U673 ( .IN1(N139), .IN2(\add_218/carry[7] ), .Q(\add_218/carry[8] ) );
  XNOR2X1 U674 ( .IN1(\add_218/carry[7] ), .IN2(N139), .Q(N537) );
  OR2X1 U675 ( .IN1(besthop[5]), .IN2(\r212/carry[6] ), .Q(\r212/carry[7] ) );
  XNOR2X1 U676 ( .IN1(\r212/carry[6] ), .IN2(besthop[5]), .Q(N168) );
  OR2X1 U677 ( .IN1(N313), .IN2(\add_151/carry[6] ), .Q(\add_151/carry[7] ) );
  XNOR2X1 U678 ( .IN1(\add_151/carry[6] ), .IN2(N313), .Q(N324) );
  AND2X1 U679 ( .IN1(\add_212/carry[6] ), .IN2(N489), .Q(\add_212/carry[7] )
         );
  XOR2X1 U680 ( .IN1(N489), .IN2(\add_212/carry[6] ), .Q(N506) );
  OR2X1 U681 ( .IN1(i[5]), .IN2(\add_137/carry[6] ), .Q(\add_137/carry[7] ) );
  XNOR2X1 U682 ( .IN1(\add_137/carry[6] ), .IN2(i[5]), .Q(N269) );
  OR2X1 U683 ( .IN1(N138), .IN2(\add_108/carry[6] ), .Q(\add_108/carry[7] ) );
  XNOR2X1 U684 ( .IN1(\add_108/carry[6] ), .IN2(N138), .Q(N155) );
  OR2X1 U685 ( .IN1(N1270), .IN2(\add_177/carry[6] ), .Q(\add_177/carry[7] )
         );
  XNOR2X1 U686 ( .IN1(\add_177/carry[6] ), .IN2(N1270), .Q(N423) );
  OR2X1 U687 ( .IN1(N138), .IN2(\add_128/carry[6] ), .Q(\add_128/carry[7] ) );
  XNOR2X1 U688 ( .IN1(\add_128/carry[6] ), .IN2(N138), .Q(N233) );
  AND2X1 U689 ( .IN1(\add_199/carry[6] ), .IN2(j[5]), .Q(\add_199/carry[7] )
         );
  XOR2X1 U690 ( .IN1(j[5]), .IN2(\add_199/carry[6] ), .Q(N477) );
  OR2X1 U691 ( .IN1(N138), .IN2(\add_218/carry[6] ), .Q(\add_218/carry[7] ) );
  XNOR2X1 U692 ( .IN1(\add_218/carry[6] ), .IN2(N138), .Q(N536) );
  OR2X1 U693 ( .IN1(i[5]), .IN2(\add_117/carry[6] ), .Q(\add_117/carry[7] ) );
  XNOR2X1 U694 ( .IN1(\add_117/carry[6] ), .IN2(i[5]), .Q(N190) );
  OR2X1 U695 ( .IN1(i[5]), .IN2(\r221/carry[6] ), .Q(\r221/carry[7] ) );
  XNOR2X1 U696 ( .IN1(\r221/carry[6] ), .IN2(i[5]), .Q(N335) );
  AND2X1 U697 ( .IN1(\add_117/carry[5] ), .IN2(i[4]), .Q(\add_117/carry[6] )
         );
  XOR2X1 U698 ( .IN1(i[4]), .IN2(\add_117/carry[5] ), .Q(N189) );
  AND2X1 U699 ( .IN1(\add_212/carry[5] ), .IN2(N488), .Q(\add_212/carry[6] )
         );
  XOR2X1 U700 ( .IN1(N488), .IN2(\add_212/carry[5] ), .Q(N505) );
  AND2X1 U701 ( .IN1(\r212/carry[5] ), .IN2(besthop[4]), .Q(\r212/carry[6] )
         );
  XOR2X1 U702 ( .IN1(besthop[4]), .IN2(\r212/carry[5] ), .Q(N167) );
  OR2X1 U703 ( .IN1(N312), .IN2(\add_151/carry[5] ), .Q(\add_151/carry[6] ) );
  XNOR2X1 U704 ( .IN1(\add_151/carry[5] ), .IN2(N312), .Q(N323) );
  AND2X1 U705 ( .IN1(\add_108/carry[5] ), .IN2(N137), .Q(\add_108/carry[6] )
         );
  XOR2X1 U706 ( .IN1(N137), .IN2(\add_108/carry[5] ), .Q(N154) );
  AND2X1 U707 ( .IN1(\add_137/carry[5] ), .IN2(i[4]), .Q(\add_137/carry[6] )
         );
  XOR2X1 U708 ( .IN1(i[4]), .IN2(\add_137/carry[5] ), .Q(N268) );
  AND2X1 U709 ( .IN1(\add_199/carry[5] ), .IN2(j[4]), .Q(\add_199/carry[6] )
         );
  XOR2X1 U710 ( .IN1(j[4]), .IN2(\add_199/carry[5] ), .Q(N476) );
  AND2X1 U711 ( .IN1(\add_177/carry[5] ), .IN2(N1272), .Q(\add_177/carry[6] )
         );
  XOR2X1 U712 ( .IN1(N1272), .IN2(\add_177/carry[5] ), .Q(N422) );
  AND2X1 U713 ( .IN1(\add_128/carry[5] ), .IN2(N137), .Q(\add_128/carry[6] )
         );
  XOR2X1 U714 ( .IN1(N137), .IN2(\add_128/carry[5] ), .Q(N232) );
  AND2X1 U715 ( .IN1(\r221/carry[5] ), .IN2(i[4]), .Q(\r221/carry[6] ) );
  XOR2X1 U716 ( .IN1(i[4]), .IN2(\r221/carry[5] ), .Q(N334) );
  AND2X1 U717 ( .IN1(\add_218/carry[5] ), .IN2(N137), .Q(\add_218/carry[6] )
         );
  XOR2X1 U718 ( .IN1(N137), .IN2(\add_218/carry[5] ), .Q(N535) );
  AND2X1 U719 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_117/carry[5] ) );
  XOR2X1 U720 ( .IN1(i[3]), .IN2(i[2]), .Q(N188) );
  AND2X1 U721 ( .IN1(N486), .IN2(N487), .Q(\add_212/carry[5] ) );
  XOR2X1 U722 ( .IN1(N487), .IN2(N486), .Q(N504) );
  AND2X1 U723 ( .IN1(besthop[2]), .IN2(besthop[3]), .Q(\r212/carry[5] ) );
  XOR2X1 U724 ( .IN1(besthop[3]), .IN2(besthop[2]), .Q(N166) );
  AND2X1 U725 ( .IN1(N310), .IN2(N311), .Q(\add_151/carry[5] ) );
  XOR2X1 U726 ( .IN1(N311), .IN2(N310), .Q(N322) );
  AND2X1 U727 ( .IN1(N135), .IN2(N136), .Q(\add_108/carry[5] ) );
  XOR2X1 U728 ( .IN1(N136), .IN2(N135), .Q(N153) );
  AND2X1 U729 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_137/carry[5] ) );
  XOR2X1 U730 ( .IN1(i[3]), .IN2(i[2]), .Q(N267) );
  AND2X1 U731 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_199/carry[5] ) );
  XOR2X1 U732 ( .IN1(j[3]), .IN2(j[2]), .Q(N475) );
  AND2X1 U733 ( .IN1(N1276), .IN2(N413), .Q(\add_177/carry[5] ) );
  XOR2X1 U734 ( .IN1(N413), .IN2(N1276), .Q(N421) );
  AND2X1 U735 ( .IN1(N135), .IN2(N136), .Q(\add_128/carry[5] ) );
  XOR2X1 U736 ( .IN1(N136), .IN2(N135), .Q(N231) );
  AND2X1 U737 ( .IN1(i[2]), .IN2(i[3]), .Q(\r221/carry[5] ) );
  XOR2X1 U738 ( .IN1(i[3]), .IN2(i[2]), .Q(N333) );
  AND2X1 U739 ( .IN1(N135), .IN2(N136), .Q(\add_218/carry[5] ) );
  XOR2X1 U740 ( .IN1(N136), .IN2(N135), .Q(N534) );
  NOR2X0 U741 ( .IN1(N293), .IN2(N292), .QN(n536) );
  AO21X1 U742 ( .IN1(N293), .IN2(N292), .IN3(n536), .Q(N320) );
  NOR2X0 U743 ( .IN1(n544), .IN2(N294), .QN(n537) );
  AO21X1 U744 ( .IN1(N294), .IN2(n544), .IN3(n537), .Q(N310) );
  NOR2X0 U745 ( .IN1(n545), .IN2(N295), .QN(n538) );
  AO21X1 U746 ( .IN1(N295), .IN2(n545), .IN3(n538), .Q(N311) );
  NOR2X0 U747 ( .IN1(n546), .IN2(N296), .QN(n539) );
  AO21X1 U748 ( .IN1(N296), .IN2(n546), .IN3(n539), .Q(N312) );
  NOR2X0 U749 ( .IN1(n547), .IN2(N297), .QN(n540) );
  AO21X1 U750 ( .IN1(N297), .IN2(n547), .IN3(n540), .Q(N313) );
  NOR2X0 U751 ( .IN1(n548), .IN2(N298), .QN(n541) );
  AO21X1 U752 ( .IN1(N298), .IN2(n548), .IN3(n541), .Q(N314) );
  NOR2X0 U753 ( .IN1(n549), .IN2(N299), .QN(n542) );
  AO21X1 U754 ( .IN1(N299), .IN2(n549), .IN3(n542), .Q(N315) );
  XNOR2X1 U755 ( .IN1(N300), .IN2(n550), .Q(N316) );
  NOR2X0 U756 ( .IN1(N300), .IN2(n550), .QN(n543) );
  XOR2X1 U757 ( .IN1(N301), .IN2(n543), .Q(N317) );
  XOR2X1 U758 ( .IN1(data_in[12]), .IN2(MY_CLUSTER_ID[12]), .Q(n554) );
  XOR2X1 U759 ( .IN1(data_in[13]), .IN2(MY_CLUSTER_ID[13]), .Q(n553) );
  XOR2X1 U760 ( .IN1(data_in[14]), .IN2(MY_CLUSTER_ID[14]), .Q(n552) );
  XOR2X1 U761 ( .IN1(data_in[15]), .IN2(MY_CLUSTER_ID[15]), .Q(n551) );
  NOR4X0 U762 ( .IN1(n554), .IN2(n553), .IN3(n552), .IN4(n551), .QN(n572) );
  XOR2X1 U763 ( .IN1(data_in[8]), .IN2(MY_CLUSTER_ID[8]), .Q(n558) );
  XOR2X1 U764 ( .IN1(data_in[9]), .IN2(MY_CLUSTER_ID[9]), .Q(n557) );
  XOR2X1 U765 ( .IN1(data_in[10]), .IN2(MY_CLUSTER_ID[10]), .Q(n556) );
  XOR2X1 U766 ( .IN1(data_in[11]), .IN2(MY_CLUSTER_ID[11]), .Q(n555) );
  NOR4X0 U767 ( .IN1(n558), .IN2(n557), .IN3(n556), .IN4(n555), .QN(n571) );
  XOR2X1 U768 ( .IN1(data_in[4]), .IN2(MY_CLUSTER_ID[4]), .Q(n562) );
  XOR2X1 U769 ( .IN1(data_in[5]), .IN2(MY_CLUSTER_ID[5]), .Q(n561) );
  XOR2X1 U770 ( .IN1(data_in[6]), .IN2(MY_CLUSTER_ID[6]), .Q(n560) );
  XOR2X1 U771 ( .IN1(data_in[7]), .IN2(MY_CLUSTER_ID[7]), .Q(n559) );
  NOR4X0 U772 ( .IN1(n562), .IN2(n561), .IN3(n560), .IN4(n559), .QN(n570) );
  NOR2X0 U773 ( .IN1(n573), .IN2(data_in[0]), .QN(n563) );
  OA22X1 U774 ( .IN1(n563), .IN2(n932), .IN3(MY_CLUSTER_ID[1]), .IN4(n563), 
        .Q(n568) );
  AND2X1 U775 ( .IN1(data_in[0]), .IN2(n573), .Q(n564) );
  OA22X1 U776 ( .IN1(data_in[1]), .IN2(n564), .IN3(n564), .IN4(n574), .Q(n567)
         );
  XOR2X1 U777 ( .IN1(data_in[2]), .IN2(MY_CLUSTER_ID[2]), .Q(n566) );
  XOR2X1 U778 ( .IN1(data_in[3]), .IN2(MY_CLUSTER_ID[3]), .Q(n565) );
  NOR4X0 U779 ( .IN1(n568), .IN2(n567), .IN3(n566), .IN4(n565), .QN(n569) );
  NAND4X0 U780 ( .IN1(n572), .IN2(n571), .IN3(n570), .IN4(n569), .QN(N130) );
  XOR2X1 U781 ( .IN1(knownSinkCount[15]), .IN2(N499), .Q(n580) );
  XOR2X1 U782 ( .IN1(knownSinkCount[2]), .IN2(N486), .Q(n579) );
  NOR2X0 U783 ( .IN1(n598), .IN2(N501), .QN(n575) );
  OA22X1 U784 ( .IN1(knownSinkCount[1]), .IN2(n575), .IN3(n575), .IN4(n597), 
        .Q(n578) );
  AND2X1 U785 ( .IN1(N501), .IN2(n598), .Q(n576) );
  OA22X1 U786 ( .IN1(n576), .IN2(n599), .IN3(N502), .IN4(n576), .Q(n577) );
  OR4X1 U787 ( .IN1(n580), .IN2(n579), .IN3(n578), .IN4(n577), .Q(n596) );
  XNOR2X1 U788 ( .IN1(knownSinkCount[6]), .IN2(N490), .Q(n584) );
  XNOR2X1 U789 ( .IN1(knownSinkCount[5]), .IN2(N489), .Q(n583) );
  XNOR2X1 U790 ( .IN1(knownSinkCount[4]), .IN2(N488), .Q(n582) );
  XNOR2X1 U791 ( .IN1(knownSinkCount[3]), .IN2(N487), .Q(n581) );
  NAND4X0 U792 ( .IN1(n584), .IN2(n583), .IN3(n582), .IN4(n581), .QN(n595) );
  XNOR2X1 U793 ( .IN1(knownSinkCount[10]), .IN2(N494), .Q(n588) );
  XNOR2X1 U794 ( .IN1(knownSinkCount[9]), .IN2(N493), .Q(n587) );
  XNOR2X1 U795 ( .IN1(knownSinkCount[8]), .IN2(N492), .Q(n586) );
  XNOR2X1 U796 ( .IN1(knownSinkCount[7]), .IN2(N491), .Q(n585) );
  NAND4X0 U797 ( .IN1(n588), .IN2(n587), .IN3(n586), .IN4(n585), .QN(n594) );
  XNOR2X1 U798 ( .IN1(knownSinkCount[14]), .IN2(N498), .Q(n592) );
  XNOR2X1 U799 ( .IN1(knownSinkCount[13]), .IN2(N497), .Q(n591) );
  XNOR2X1 U800 ( .IN1(knownSinkCount[12]), .IN2(N496), .Q(n590) );
  XNOR2X1 U801 ( .IN1(knownSinkCount[11]), .IN2(N495), .Q(n589) );
  NAND4X0 U802 ( .IN1(n592), .IN2(n591), .IN3(n590), .IN4(n589), .QN(n593) );
  NOR4X0 U803 ( .IN1(n596), .IN2(n595), .IN3(n594), .IN4(n593), .QN(N511) );
  XOR2X1 U804 ( .IN1(neighborCount[15]), .IN2(N148), .Q(n605) );
  XOR2X1 U805 ( .IN1(neighborCount[2]), .IN2(N135), .Q(n604) );
  NOR2X0 U806 ( .IN1(n624), .IN2(N150), .QN(n600) );
  OA22X1 U807 ( .IN1(neighborCount[1]), .IN2(n600), .IN3(n600), .IN4(n623), 
        .Q(n603) );
  AND2X1 U808 ( .IN1(N150), .IN2(n624), .Q(n601) );
  OA22X1 U809 ( .IN1(n601), .IN2(n622), .IN3(N151), .IN4(n601), .Q(n602) );
  OR4X1 U810 ( .IN1(n605), .IN2(n604), .IN3(n603), .IN4(n602), .Q(n621) );
  XNOR2X1 U811 ( .IN1(neighborCount[6]), .IN2(N139), .Q(n609) );
  XNOR2X1 U812 ( .IN1(neighborCount[5]), .IN2(N138), .Q(n608) );
  XNOR2X1 U813 ( .IN1(neighborCount[4]), .IN2(N137), .Q(n607) );
  XNOR2X1 U814 ( .IN1(neighborCount[3]), .IN2(N136), .Q(n606) );
  NAND4X0 U815 ( .IN1(n609), .IN2(n608), .IN3(n607), .IN4(n606), .QN(n620) );
  XNOR2X1 U816 ( .IN1(neighborCount[10]), .IN2(N143), .Q(n613) );
  XNOR2X1 U817 ( .IN1(neighborCount[9]), .IN2(N142), .Q(n612) );
  XNOR2X1 U818 ( .IN1(neighborCount[8]), .IN2(N141), .Q(n611) );
  XNOR2X1 U819 ( .IN1(neighborCount[7]), .IN2(N140), .Q(n610) );
  NAND4X0 U820 ( .IN1(n613), .IN2(n612), .IN3(n611), .IN4(n610), .QN(n619) );
  XNOR2X1 U821 ( .IN1(neighborCount[14]), .IN2(N147), .Q(n617) );
  XNOR2X1 U822 ( .IN1(neighborCount[13]), .IN2(N146), .Q(n616) );
  XNOR2X1 U823 ( .IN1(neighborCount[12]), .IN2(N145), .Q(n615) );
  XNOR2X1 U824 ( .IN1(neighborCount[11]), .IN2(N144), .Q(n614) );
  NAND4X0 U825 ( .IN1(n617), .IN2(n616), .IN3(n615), .IN4(n614), .QN(n618) );
  NOR4X0 U826 ( .IN1(n621), .IN2(n620), .IN3(n619), .IN4(n618), .QN(N160) );
  NOR2X0 U827 ( .IN1(k[11]), .IN2(k[10]), .QN(n630) );
  AO21X1 U828 ( .IN1(k[1]), .IN2(k[0]), .IN3(k[2]), .Q(n625) );
  NAND2X0 U829 ( .IN1(k[3]), .IN2(n625), .QN(n629) );
  NOR3X0 U830 ( .IN1(k[12]), .IN2(k[14]), .IN3(k[13]), .QN(n628) );
  OR4X1 U831 ( .IN1(k[7]), .IN2(k[6]), .IN3(k[9]), .IN4(k[8]), .Q(n626) );
  NOR4X0 U832 ( .IN1(n626), .IN2(k[15]), .IN3(k[5]), .IN4(k[4]), .QN(n627) );
  NAND4X0 U833 ( .IN1(n630), .IN2(n629), .IN3(n628), .IN4(n627), .QN(N406) );
  AND2X1 U834 ( .IN1(n662), .IN2(bestvalue[14]), .Q(n646) );
  NOR2X0 U835 ( .IN1(n648), .IN2(N441), .QN(n631) );
  AND2X1 U836 ( .IN1(n649), .IN2(n631), .Q(n632) );
  OA222X1 U837 ( .IN1(bestvalue[2]), .IN2(n650), .IN3(bestvalue[1]), .IN4(n632), .IN5(n631), .IN6(n649), .Q(n633) );
  AO221X1 U838 ( .IN1(bestvalue[2]), .IN2(n650), .IN3(bestvalue[3]), .IN4(n651), .IN5(n633), .Q(n634) );
  OA221X1 U839 ( .IN1(bestvalue[4]), .IN2(n652), .IN3(bestvalue[3]), .IN4(n651), .IN5(n634), .Q(n635) );
  AO221X1 U840 ( .IN1(bestvalue[4]), .IN2(n652), .IN3(bestvalue[5]), .IN4(n653), .IN5(n635), .Q(n636) );
  OA221X1 U841 ( .IN1(bestvalue[6]), .IN2(n654), .IN3(bestvalue[5]), .IN4(n653), .IN5(n636), .Q(n637) );
  AO221X1 U842 ( .IN1(bestvalue[6]), .IN2(n654), .IN3(bestvalue[7]), .IN4(n655), .IN5(n637), .Q(n638) );
  OA221X1 U843 ( .IN1(bestvalue[8]), .IN2(n656), .IN3(bestvalue[7]), .IN4(n655), .IN5(n638), .Q(n639) );
  AO221X1 U844 ( .IN1(bestvalue[8]), .IN2(n656), .IN3(bestvalue[9]), .IN4(n657), .IN5(n639), .Q(n640) );
  OA221X1 U845 ( .IN1(bestvalue[9]), .IN2(n657), .IN3(bestvalue[10]), .IN4(
        n658), .IN5(n640), .Q(n641) );
  AO221X1 U846 ( .IN1(bestvalue[10]), .IN2(n658), .IN3(bestvalue[11]), .IN4(
        n659), .IN5(n641), .Q(n642) );
  OA221X1 U847 ( .IN1(bestvalue[12]), .IN2(n660), .IN3(bestvalue[11]), .IN4(
        n659), .IN5(n642), .Q(n643) );
  AO221X1 U848 ( .IN1(bestvalue[12]), .IN2(n660), .IN3(bestvalue[13]), .IN4(
        n661), .IN5(n643), .Q(n644) );
  OA221X1 U849 ( .IN1(bestvalue[14]), .IN2(n662), .IN3(bestvalue[13]), .IN4(
        n661), .IN5(n644), .Q(n645) );
  OA22X1 U850 ( .IN1(bestvalue[15]), .IN2(n663), .IN3(n646), .IN4(n645), .Q(
        n647) );
  AO21X1 U851 ( .IN1(bestvalue[15]), .IN2(n663), .IN3(n647), .Q(N459) );
  XOR2X1 U852 ( .IN1(data_in[15]), .IN2(neighborID[15]), .Q(n669) );
  XOR2X1 U853 ( .IN1(data_in[2]), .IN2(neighborID[2]), .Q(n668) );
  NOR2X0 U854 ( .IN1(n933), .IN2(neighborID[0]), .QN(n664) );
  OA22X1 U855 ( .IN1(data_in[1]), .IN2(n664), .IN3(n664), .IN4(n686), .Q(n667)
         );
  AND2X1 U856 ( .IN1(neighborID[0]), .IN2(n933), .Q(n665) );
  OA22X1 U857 ( .IN1(n665), .IN2(n932), .IN3(neighborID[1]), .IN4(n665), .Q(
        n666) );
  OR4X1 U858 ( .IN1(n669), .IN2(n668), .IN3(n667), .IN4(n666), .Q(n685) );
  XNOR2X1 U859 ( .IN1(data_in[6]), .IN2(neighborID[6]), .Q(n673) );
  XNOR2X1 U860 ( .IN1(data_in[5]), .IN2(neighborID[5]), .Q(n672) );
  XNOR2X1 U861 ( .IN1(data_in[4]), .IN2(neighborID[4]), .Q(n671) );
  XNOR2X1 U862 ( .IN1(data_in[3]), .IN2(neighborID[3]), .Q(n670) );
  NAND4X0 U863 ( .IN1(n673), .IN2(n672), .IN3(n671), .IN4(n670), .QN(n684) );
  XNOR2X1 U864 ( .IN1(data_in[10]), .IN2(neighborID[10]), .Q(n677) );
  XNOR2X1 U865 ( .IN1(data_in[9]), .IN2(neighborID[9]), .Q(n676) );
  XNOR2X1 U866 ( .IN1(data_in[8]), .IN2(neighborID[8]), .Q(n675) );
  XNOR2X1 U867 ( .IN1(data_in[7]), .IN2(neighborID[7]), .Q(n674) );
  NAND4X0 U868 ( .IN1(n677), .IN2(n676), .IN3(n675), .IN4(n674), .QN(n683) );
  XNOR2X1 U869 ( .IN1(data_in[14]), .IN2(neighborID[14]), .Q(n681) );
  XNOR2X1 U870 ( .IN1(data_in[13]), .IN2(neighborID[13]), .Q(n680) );
  XNOR2X1 U871 ( .IN1(data_in[12]), .IN2(neighborID[12]), .Q(n679) );
  XNOR2X1 U872 ( .IN1(data_in[11]), .IN2(neighborID[11]), .Q(n678) );
  NAND4X0 U873 ( .IN1(n681), .IN2(n680), .IN3(n679), .IN4(n678), .QN(n682) );
  NOR4X0 U874 ( .IN1(n685), .IN2(n684), .IN3(n683), .IN4(n682), .QN(N483) );
  AO22X1 U875 ( .IN1(n687), .IN2(neighborCount[0]), .IN3(data_in[0]), .IN4(
        n688), .Q(n527) );
  MUX21X1 U876 ( .IN1(n689), .IN2(state[3]), .S(n690), .Q(n526) );
  NAND4X0 U877 ( .IN1(n691), .IN2(n692), .IN3(n693), .IN4(n694), .QN(n689) );
  AND4X1 U878 ( .IN1(n695), .IN2(n696), .IN3(n697), .IN4(n698), .Q(n694) );
  OA21X1 U879 ( .IN1(n699), .IN2(n700), .IN3(nrst), .Q(n693) );
  NAND4X0 U880 ( .IN1(n701), .IN2(n702), .IN3(n703), .IN4(n704), .QN(n525) );
  NOR2X0 U881 ( .IN1(n705), .IN2(n706), .QN(n704) );
  NAND2X0 U882 ( .IN1(n707), .IN2(n699), .QN(n703) );
  NAND4X0 U883 ( .IN1(n708), .IN2(n709), .IN3(n701), .IN4(n710), .QN(n524) );
  NOR2X0 U884 ( .IN1(n711), .IN2(n705), .QN(n710) );
  NAND3X0 U885 ( .IN1(n712), .IN2(nrst), .IN3(n713), .QN(n705) );
  OA22X1 U886 ( .IN1(N160), .IN2(n714), .IN3(en), .IN4(n715), .Q(n713) );
  NOR2X0 U887 ( .IN1(n690), .IN2(n716), .QN(n523) );
  NOR4X0 U888 ( .IN1(n717), .IN2(n718), .IN3(n719), .IN4(n720), .QN(n716) );
  INVX0 U889 ( .INP(n692), .ZN(n720) );
  OA221X1 U890 ( .IN1(n699), .IN2(n714), .IN3(n715), .IN4(en), .IN5(n721), .Q(
        n692) );
  AND2X1 U891 ( .IN1(n722), .IN2(n723), .Q(n721) );
  NOR2X0 U892 ( .IN1(n699), .IN2(n724), .QN(n719) );
  NAND3X0 U893 ( .IN1(n725), .IN2(n702), .IN3(n726), .QN(n717) );
  INVX0 U894 ( .INP(n701), .ZN(n690) );
  NAND4X0 U895 ( .IN1(n727), .IN2(n697), .IN3(n728), .IN4(n729), .QN(n701) );
  NOR4X0 U896 ( .IN1(n730), .IN2(n711), .IN3(n731), .IN4(n732), .QN(n729) );
  NOR2X0 U897 ( .IN1(n699), .IN2(n725), .QN(n732) );
  INVX0 U898 ( .INP(n712), .ZN(n731) );
  NOR2X0 U899 ( .IN1(n733), .IN2(n734), .QN(n712) );
  NAND3X0 U900 ( .IN1(n735), .IN2(n736), .IN3(n723), .QN(n711) );
  NOR3X0 U901 ( .IN1(n707), .IN2(n737), .IN3(n738), .QN(n728) );
  AO22X1 U902 ( .IN1(n739), .IN2(batteryStat[0]), .IN3(n740), .IN4(data_in[0]), 
        .Q(n522) );
  AO22X1 U903 ( .IN1(n739), .IN2(batteryStat[1]), .IN3(n740), .IN4(data_in[1]), 
        .Q(n521) );
  AO22X1 U904 ( .IN1(n739), .IN2(batteryStat[2]), .IN3(n740), .IN4(data_in[2]), 
        .Q(n520) );
  AO22X1 U905 ( .IN1(n739), .IN2(batteryStat[3]), .IN3(n740), .IN4(data_in[3]), 
        .Q(n519) );
  AO22X1 U906 ( .IN1(n739), .IN2(batteryStat[4]), .IN3(n740), .IN4(data_in[4]), 
        .Q(n518) );
  AO22X1 U907 ( .IN1(n739), .IN2(batteryStat[5]), .IN3(n740), .IN4(data_in[5]), 
        .Q(n517) );
  AO22X1 U908 ( .IN1(n739), .IN2(batteryStat[6]), .IN3(n740), .IN4(data_in[6]), 
        .Q(n516) );
  AO22X1 U909 ( .IN1(n739), .IN2(batteryStat[7]), .IN3(n740), .IN4(data_in[7]), 
        .Q(n515) );
  AO22X1 U910 ( .IN1(n739), .IN2(batteryStat[8]), .IN3(n740), .IN4(data_in[8]), 
        .Q(n514) );
  AO22X1 U911 ( .IN1(n739), .IN2(batteryStat[9]), .IN3(n740), .IN4(data_in[9]), 
        .Q(n513) );
  AO22X1 U912 ( .IN1(n739), .IN2(batteryStat[10]), .IN3(n740), .IN4(
        data_in[10]), .Q(n512) );
  AO22X1 U913 ( .IN1(n739), .IN2(batteryStat[11]), .IN3(n740), .IN4(
        data_in[11]), .Q(n511) );
  AO22X1 U914 ( .IN1(n739), .IN2(batteryStat[12]), .IN3(n740), .IN4(
        data_in[12]), .Q(n510) );
  AO22X1 U915 ( .IN1(n739), .IN2(batteryStat[13]), .IN3(n740), .IN4(
        data_in[13]), .Q(n509) );
  AO22X1 U916 ( .IN1(n739), .IN2(batteryStat[14]), .IN3(n740), .IN4(
        data_in[14]), .Q(n508) );
  AO22X1 U917 ( .IN1(n739), .IN2(batteryStat[15]), .IN3(n740), .IN4(
        data_in[15]), .Q(n507) );
  AO22X1 U918 ( .IN1(n743), .IN2(neighborID[0]), .IN3(n744), .IN4(data_in[0]), 
        .Q(n506) );
  AO22X1 U919 ( .IN1(n743), .IN2(neighborID[1]), .IN3(n744), .IN4(data_in[1]), 
        .Q(n505) );
  AO22X1 U920 ( .IN1(n743), .IN2(neighborID[2]), .IN3(n744), .IN4(data_in[2]), 
        .Q(n504) );
  AO22X1 U921 ( .IN1(n743), .IN2(neighborID[3]), .IN3(n744), .IN4(data_in[3]), 
        .Q(n503) );
  AO22X1 U922 ( .IN1(n743), .IN2(neighborID[4]), .IN3(n744), .IN4(data_in[4]), 
        .Q(n502) );
  AO22X1 U923 ( .IN1(n743), .IN2(neighborID[5]), .IN3(n744), .IN4(data_in[5]), 
        .Q(n501) );
  AO22X1 U924 ( .IN1(n743), .IN2(neighborID[6]), .IN3(n744), .IN4(data_in[6]), 
        .Q(n500) );
  AO22X1 U925 ( .IN1(n743), .IN2(neighborID[7]), .IN3(n744), .IN4(data_in[7]), 
        .Q(n499) );
  AO22X1 U926 ( .IN1(n743), .IN2(neighborID[8]), .IN3(n744), .IN4(data_in[8]), 
        .Q(n498) );
  AO22X1 U927 ( .IN1(n743), .IN2(neighborID[9]), .IN3(n744), .IN4(data_in[9]), 
        .Q(n497) );
  AO22X1 U928 ( .IN1(n743), .IN2(neighborID[10]), .IN3(n744), .IN4(data_in[10]), .Q(n496) );
  AO22X1 U929 ( .IN1(n743), .IN2(neighborID[11]), .IN3(n744), .IN4(data_in[11]), .Q(n495) );
  AO22X1 U930 ( .IN1(n743), .IN2(neighborID[12]), .IN3(n744), .IN4(data_in[12]), .Q(n494) );
  AO22X1 U931 ( .IN1(n743), .IN2(neighborID[13]), .IN3(n744), .IN4(data_in[13]), .Q(n493) );
  AO22X1 U932 ( .IN1(n743), .IN2(neighborID[14]), .IN3(n744), .IN4(data_in[14]), .Q(n492) );
  AO22X1 U933 ( .IN1(n743), .IN2(neighborID[15]), .IN3(n744), .IN4(data_in[15]), .Q(n491) );
  AO22X1 U934 ( .IN1(n687), .IN2(neighborCount[1]), .IN3(data_in[1]), .IN4(
        n688), .Q(n490) );
  AO22X1 U935 ( .IN1(n687), .IN2(neighborCount[2]), .IN3(data_in[2]), .IN4(
        n688), .Q(n489) );
  AO22X1 U936 ( .IN1(n687), .IN2(neighborCount[3]), .IN3(data_in[3]), .IN4(
        n688), .Q(n488) );
  AO22X1 U937 ( .IN1(n687), .IN2(neighborCount[4]), .IN3(data_in[4]), .IN4(
        n688), .Q(n487) );
  AO22X1 U938 ( .IN1(n687), .IN2(neighborCount[5]), .IN3(data_in[5]), .IN4(
        n688), .Q(n486) );
  AO22X1 U939 ( .IN1(n687), .IN2(neighborCount[6]), .IN3(data_in[6]), .IN4(
        n688), .Q(n485) );
  AO22X1 U940 ( .IN1(n687), .IN2(neighborCount[7]), .IN3(data_in[7]), .IN4(
        n688), .Q(n484) );
  AO22X1 U941 ( .IN1(n687), .IN2(neighborCount[8]), .IN3(data_in[8]), .IN4(
        n688), .Q(n483) );
  AO22X1 U942 ( .IN1(n687), .IN2(neighborCount[9]), .IN3(data_in[9]), .IN4(
        n688), .Q(n482) );
  AO22X1 U943 ( .IN1(n687), .IN2(neighborCount[10]), .IN3(data_in[10]), .IN4(
        n688), .Q(n481) );
  AO22X1 U944 ( .IN1(n687), .IN2(neighborCount[11]), .IN3(data_in[11]), .IN4(
        n688), .Q(n480) );
  AO22X1 U945 ( .IN1(n687), .IN2(neighborCount[12]), .IN3(data_in[12]), .IN4(
        n688), .Q(n479) );
  AO22X1 U946 ( .IN1(n687), .IN2(neighborCount[13]), .IN3(data_in[13]), .IN4(
        n688), .Q(n478) );
  AO22X1 U947 ( .IN1(n687), .IN2(neighborCount[14]), .IN3(data_in[14]), .IN4(
        n688), .Q(n477) );
  AO22X1 U948 ( .IN1(n687), .IN2(neighborCount[15]), .IN3(data_in[15]), .IN4(
        n688), .Q(n476) );
  AO22X1 U949 ( .IN1(n749), .IN2(knownSinkCount[0]), .IN3(n750), .IN4(
        data_in[0]), .Q(n475) );
  AO22X1 U950 ( .IN1(n749), .IN2(knownSinkCount[1]), .IN3(n750), .IN4(
        data_in[1]), .Q(n474) );
  AO22X1 U951 ( .IN1(n749), .IN2(knownSinkCount[2]), .IN3(n750), .IN4(
        data_in[2]), .Q(n473) );
  AO22X1 U952 ( .IN1(n749), .IN2(knownSinkCount[3]), .IN3(n750), .IN4(
        data_in[3]), .Q(n472) );
  AO22X1 U953 ( .IN1(n749), .IN2(knownSinkCount[4]), .IN3(n750), .IN4(
        data_in[4]), .Q(n471) );
  AO22X1 U954 ( .IN1(n749), .IN2(knownSinkCount[5]), .IN3(n750), .IN4(
        data_in[5]), .Q(n470) );
  AO22X1 U955 ( .IN1(n749), .IN2(knownSinkCount[6]), .IN3(n750), .IN4(
        data_in[6]), .Q(n469) );
  AO22X1 U956 ( .IN1(n749), .IN2(knownSinkCount[7]), .IN3(n750), .IN4(
        data_in[7]), .Q(n468) );
  AO22X1 U957 ( .IN1(n749), .IN2(knownSinkCount[8]), .IN3(n750), .IN4(
        data_in[8]), .Q(n467) );
  AO22X1 U958 ( .IN1(n749), .IN2(knownSinkCount[9]), .IN3(n750), .IN4(
        data_in[9]), .Q(n466) );
  AO22X1 U959 ( .IN1(n749), .IN2(knownSinkCount[10]), .IN3(n750), .IN4(
        data_in[10]), .Q(n465) );
  AO22X1 U960 ( .IN1(n749), .IN2(knownSinkCount[11]), .IN3(n750), .IN4(
        data_in[11]), .Q(n464) );
  AO22X1 U961 ( .IN1(n749), .IN2(knownSinkCount[12]), .IN3(n750), .IN4(
        data_in[12]), .Q(n463) );
  AO22X1 U962 ( .IN1(n749), .IN2(knownSinkCount[13]), .IN3(n750), .IN4(
        data_in[13]), .Q(n462) );
  AO22X1 U963 ( .IN1(n749), .IN2(knownSinkCount[14]), .IN3(n750), .IN4(
        data_in[14]), .Q(n461) );
  AO22X1 U964 ( .IN1(n749), .IN2(knownSinkCount[15]), .IN3(n750), .IN4(
        data_in[15]), .Q(n460) );
  AO22X1 U965 ( .IN1(n752), .IN2(N472), .IN3(N501), .IN4(n753), .Q(n459) );
  AO22X1 U966 ( .IN1(n752), .IN2(N473), .IN3(N502), .IN4(n753), .Q(n458) );
  AO22X1 U967 ( .IN1(n752), .IN2(j[2]), .IN3(N486), .IN4(n753), .Q(n457) );
  AO22X1 U968 ( .IN1(n752), .IN2(j[3]), .IN3(N487), .IN4(n753), .Q(n456) );
  AO22X1 U969 ( .IN1(n752), .IN2(j[4]), .IN3(N488), .IN4(n753), .Q(n455) );
  AO22X1 U970 ( .IN1(n752), .IN2(j[5]), .IN3(N489), .IN4(n753), .Q(n454) );
  AO22X1 U971 ( .IN1(n752), .IN2(j[6]), .IN3(N490), .IN4(n753), .Q(n453) );
  AO22X1 U972 ( .IN1(n752), .IN2(j[7]), .IN3(N491), .IN4(n753), .Q(n452) );
  AO22X1 U973 ( .IN1(n752), .IN2(j[8]), .IN3(N492), .IN4(n753), .Q(n451) );
  AO22X1 U974 ( .IN1(n752), .IN2(j[9]), .IN3(N493), .IN4(n753), .Q(n450) );
  AO22X1 U975 ( .IN1(n752), .IN2(j[10]), .IN3(N494), .IN4(n753), .Q(n449) );
  AO22X1 U976 ( .IN1(n752), .IN2(j[11]), .IN3(N495), .IN4(n753), .Q(n448) );
  AO22X1 U977 ( .IN1(n752), .IN2(j[12]), .IN3(N496), .IN4(n753), .Q(n447) );
  AO22X1 U978 ( .IN1(n752), .IN2(j[13]), .IN3(N497), .IN4(n753), .Q(n446) );
  AO22X1 U979 ( .IN1(n752), .IN2(j[14]), .IN3(N498), .IN4(n753), .Q(n445) );
  AO22X1 U980 ( .IN1(n752), .IN2(j[15]), .IN3(N499), .IN4(n753), .Q(n444) );
  AO22X1 U981 ( .IN1(n756), .IN2(i[15]), .IN3(N148), .IN4(n757), .Q(n443) );
  AO22X1 U982 ( .IN1(n756), .IN2(N330), .IN3(N150), .IN4(n757), .Q(n442) );
  AO22X1 U983 ( .IN1(n756), .IN2(N331), .IN3(N151), .IN4(n757), .Q(n441) );
  AO22X1 U984 ( .IN1(n756), .IN2(i[2]), .IN3(N135), .IN4(n757), .Q(n440) );
  AO22X1 U985 ( .IN1(n756), .IN2(i[3]), .IN3(N136), .IN4(n757), .Q(n439) );
  AO22X1 U986 ( .IN1(n756), .IN2(i[4]), .IN3(N137), .IN4(n757), .Q(n438) );
  AO22X1 U987 ( .IN1(n756), .IN2(i[5]), .IN3(N138), .IN4(n757), .Q(n437) );
  AO22X1 U988 ( .IN1(n756), .IN2(i[6]), .IN3(N139), .IN4(n757), .Q(n436) );
  AO22X1 U989 ( .IN1(n756), .IN2(i[7]), .IN3(N140), .IN4(n757), .Q(n435) );
  AO22X1 U990 ( .IN1(n756), .IN2(i[8]), .IN3(N141), .IN4(n757), .Q(n434) );
  AO22X1 U991 ( .IN1(n756), .IN2(i[9]), .IN3(N142), .IN4(n757), .Q(n433) );
  AO22X1 U992 ( .IN1(n756), .IN2(i[10]), .IN3(N143), .IN4(n757), .Q(n432) );
  AO22X1 U993 ( .IN1(n756), .IN2(i[11]), .IN3(N144), .IN4(n757), .Q(n431) );
  AO22X1 U994 ( .IN1(n756), .IN2(i[12]), .IN3(N145), .IN4(n757), .Q(n430) );
  AO22X1 U995 ( .IN1(n756), .IN2(i[13]), .IN3(N146), .IN4(n757), .Q(n429) );
  AO22X1 U996 ( .IN1(n756), .IN2(i[14]), .IN3(N147), .IN4(n757), .Q(n428) );
  AO21X1 U997 ( .IN1(n760), .IN2(N330), .IN3(n761), .Q(n427) );
  MUX21X1 U998 ( .IN1(nextsinks[0]), .IN2(n762), .S(n763), .Q(n761) );
  AO22X1 U999 ( .IN1(nextsinks[1]), .IN2(n764), .IN3(n765), .IN4(N331), .Q(
        n426) );
  AO22X1 U1000 ( .IN1(nextsinks[2]), .IN2(n764), .IN3(n765), .IN4(i[2]), .Q(
        n425) );
  AO22X1 U1001 ( .IN1(nextsinks[3]), .IN2(n764), .IN3(n765), .IN4(i[3]), .Q(
        n424) );
  AO22X1 U1002 ( .IN1(nextsinks[4]), .IN2(n764), .IN3(n765), .IN4(i[4]), .Q(
        n423) );
  AO22X1 U1003 ( .IN1(nextsinks[5]), .IN2(n764), .IN3(n765), .IN4(i[5]), .Q(
        n422) );
  AO21X1 U1004 ( .IN1(n760), .IN2(i[6]), .IN3(n766), .Q(n421) );
  MUX21X1 U1005 ( .IN1(nextsinks[6]), .IN2(n762), .S(n763), .Q(n766) );
  AO22X1 U1006 ( .IN1(nextsinks[7]), .IN2(n764), .IN3(n765), .IN4(i[7]), .Q(
        n420) );
  AO22X1 U1007 ( .IN1(nextsinks[8]), .IN2(n764), .IN3(n765), .IN4(i[8]), .Q(
        n419) );
  AO22X1 U1008 ( .IN1(nextsinks[9]), .IN2(n764), .IN3(n765), .IN4(i[9]), .Q(
        n418) );
  AO22X1 U1009 ( .IN1(nextsinks[10]), .IN2(n764), .IN3(n765), .IN4(i[10]), .Q(
        n417) );
  AO22X1 U1010 ( .IN1(nextsinks[11]), .IN2(n764), .IN3(n765), .IN4(i[11]), .Q(
        n416) );
  AO22X1 U1011 ( .IN1(nextsinks[12]), .IN2(n764), .IN3(n765), .IN4(i[12]), .Q(
        n415) );
  AO22X1 U1012 ( .IN1(nextsinks[13]), .IN2(n764), .IN3(n765), .IN4(i[13]), .Q(
        n414) );
  AO22X1 U1013 ( .IN1(nextsinks[14]), .IN2(n764), .IN3(n765), .IN4(i[14]), .Q(
        n413) );
  AO22X1 U1014 ( .IN1(nextsinks[15]), .IN2(n764), .IN3(n765), .IN4(i[15]), .Q(
        n412) );
  NOR2X0 U1015 ( .IN1(n714), .IN2(n764), .QN(n760) );
  AO21X1 U1016 ( .IN1(N483), .IN2(n755), .IN3(n742), .Q(n763) );
  AO22X1 U1017 ( .IN1(N458), .IN2(n533), .IN3(n534), .IN4(fpTemp[30]), .Q(n411) );
  AO22X1 U1018 ( .IN1(N457), .IN2(n533), .IN3(n534), .IN4(fpTemp[29]), .Q(n410) );
  AO22X1 U1019 ( .IN1(N456), .IN2(n533), .IN3(n534), .IN4(fpTemp[28]), .Q(n409) );
  AO22X1 U1020 ( .IN1(N455), .IN2(n533), .IN3(n534), .IN4(fpTemp[27]), .Q(n408) );
  AO22X1 U1021 ( .IN1(N454), .IN2(n533), .IN3(n534), .IN4(fpTemp[26]), .Q(n407) );
  AO22X1 U1022 ( .IN1(N453), .IN2(n533), .IN3(n534), .IN4(fpTemp[25]), .Q(n406) );
  AO22X1 U1023 ( .IN1(N452), .IN2(n533), .IN3(n534), .IN4(fpTemp[24]), .Q(n405) );
  AO22X1 U1024 ( .IN1(N451), .IN2(n533), .IN3(n534), .IN4(fpTemp[23]), .Q(n404) );
  AO22X1 U1025 ( .IN1(N450), .IN2(n533), .IN3(n534), .IN4(fpTemp[22]), .Q(n403) );
  AO22X1 U1026 ( .IN1(N449), .IN2(n533), .IN3(n534), .IN4(fpTemp[21]), .Q(n402) );
  AO22X1 U1027 ( .IN1(N448), .IN2(n533), .IN3(n534), .IN4(fpTemp[20]), .Q(n401) );
  AO222X1 U1028 ( .IN1(n535), .IN2(fpTemp[19]), .IN3(N371), .IN4(n767), .IN5(
        N447), .IN6(n532), .Q(n400) );
  AO222X1 U1029 ( .IN1(n534), .IN2(fpTemp[18]), .IN3(N370), .IN4(n767), .IN5(
        N446), .IN6(n532), .Q(n399) );
  AO222X1 U1030 ( .IN1(n534), .IN2(fpTemp[17]), .IN3(N369), .IN4(n767), .IN5(
        N445), .IN6(n532), .Q(n398) );
  AO222X1 U1031 ( .IN1(n535), .IN2(fpTemp[16]), .IN3(N368), .IN4(n767), .IN5(
        N444), .IN6(n532), .Q(n397) );
  AO222X1 U1032 ( .IN1(n534), .IN2(fpTemp[15]), .IN3(N367), .IN4(n767), .IN5(
        N443), .IN6(n532), .Q(n396) );
  AO222X1 U1033 ( .IN1(n535), .IN2(n768), .IN3(N366), .IN4(n767), .IN5(N442), 
        .IN6(n532), .Q(n395) );
  AO222X1 U1034 ( .IN1(n534), .IN2(n769), .IN3(N365), .IN4(n767), .IN5(N441), 
        .IN6(n532), .Q(n394) );
  AO222X1 U1035 ( .IN1(n535), .IN2(n770), .IN3(N364), .IN4(n767), .IN5(N440), 
        .IN6(n532), .Q(n393) );
  AO222X1 U1036 ( .IN1(n535), .IN2(n771), .IN3(N363), .IN4(n767), .IN5(N439), 
        .IN6(n532), .Q(n392) );
  AO222X1 U1037 ( .IN1(n535), .IN2(n772), .IN3(N362), .IN4(n767), .IN5(N438), 
        .IN6(n532), .Q(n391) );
  AO222X1 U1038 ( .IN1(n535), .IN2(n773), .IN3(N361), .IN4(n767), .IN5(N437), 
        .IN6(n531), .Q(n390) );
  AO222X1 U1039 ( .IN1(n535), .IN2(n774), .IN3(N360), .IN4(n767), .IN5(N436), 
        .IN6(n532), .Q(n389) );
  AO222X1 U1040 ( .IN1(n535), .IN2(n775), .IN3(N359), .IN4(n767), .IN5(N435), 
        .IN6(n531), .Q(n388) );
  AO222X1 U1041 ( .IN1(n535), .IN2(n776), .IN3(N358), .IN4(n767), .IN5(N434), 
        .IN6(n531), .Q(n387) );
  AO222X1 U1042 ( .IN1(n535), .IN2(n777), .IN3(N357), .IN4(n767), .IN5(N433), 
        .IN6(n531), .Q(n386) );
  AO222X1 U1043 ( .IN1(n535), .IN2(n778), .IN3(N356), .IN4(n767), .IN5(N432), 
        .IN6(n531), .Q(n385) );
  AO222X1 U1044 ( .IN1(n535), .IN2(n779), .IN3(N355), .IN4(n767), .IN5(N431), 
        .IN6(n531), .Q(n384) );
  AO222X1 U1045 ( .IN1(n535), .IN2(n780), .IN3(N354), .IN4(n767), .IN5(N430), 
        .IN6(n531), .Q(n383) );
  AO222X1 U1046 ( .IN1(n535), .IN2(n781), .IN3(N353), .IN4(n767), .IN5(N429), 
        .IN6(n531), .Q(n382) );
  AO22X1 U1047 ( .IN1(N428), .IN2(n532), .IN3(n534), .IN4(n782), .Q(n381) );
  INVX0 U1048 ( .INP(n726), .ZN(n734) );
  AO222X1 U1049 ( .IN1(n784), .IN2(fpTemp[30]), .IN3(n785), .IN4(k[15]), .IN5(
        N389), .IN6(n786), .Q(n380) );
  AO222X1 U1050 ( .IN1(n784), .IN2(fpTemp[15]), .IN3(n785), .IN4(k[0]), .IN5(
        N374), .IN6(n786), .Q(n379) );
  AO221X1 U1051 ( .IN1(n784), .IN2(fpTemp[16]), .IN3(N375), .IN4(n786), .IN5(
        n787), .Q(n378) );
  AO21X1 U1052 ( .IN1(n785), .IN2(k[1]), .IN3(n788), .Q(n787) );
  AO222X1 U1053 ( .IN1(n784), .IN2(fpTemp[17]), .IN3(n785), .IN4(k[2]), .IN5(
        N376), .IN6(n786), .Q(n377) );
  AO221X1 U1054 ( .IN1(n784), .IN2(fpTemp[18]), .IN3(N377), .IN4(n786), .IN5(
        n789), .Q(n376) );
  AO21X1 U1055 ( .IN1(n785), .IN2(k[3]), .IN3(n788), .Q(n789) );
  NOR3X0 U1056 ( .IN1(n741), .IN2(n785), .IN3(n695), .QN(n788) );
  AO222X1 U1057 ( .IN1(n784), .IN2(fpTemp[19]), .IN3(n785), .IN4(k[4]), .IN5(
        N378), .IN6(n786), .Q(n375) );
  AO222X1 U1058 ( .IN1(n784), .IN2(fpTemp[20]), .IN3(n785), .IN4(k[5]), .IN5(
        N379), .IN6(n786), .Q(n374) );
  AO222X1 U1059 ( .IN1(n784), .IN2(fpTemp[21]), .IN3(n785), .IN4(k[6]), .IN5(
        N380), .IN6(n786), .Q(n373) );
  AO222X1 U1060 ( .IN1(n784), .IN2(fpTemp[22]), .IN3(n785), .IN4(k[7]), .IN5(
        N381), .IN6(n786), .Q(n372) );
  AO222X1 U1061 ( .IN1(n784), .IN2(fpTemp[23]), .IN3(n785), .IN4(k[8]), .IN5(
        N382), .IN6(n786), .Q(n371) );
  AO222X1 U1062 ( .IN1(n784), .IN2(fpTemp[24]), .IN3(n785), .IN4(k[9]), .IN5(
        N383), .IN6(n786), .Q(n370) );
  AO222X1 U1063 ( .IN1(n784), .IN2(fpTemp[25]), .IN3(n785), .IN4(k[10]), .IN5(
        N384), .IN6(n786), .Q(n369) );
  AO222X1 U1064 ( .IN1(n784), .IN2(fpTemp[26]), .IN3(n785), .IN4(k[11]), .IN5(
        N385), .IN6(n786), .Q(n368) );
  AO222X1 U1065 ( .IN1(n784), .IN2(fpTemp[27]), .IN3(n785), .IN4(k[12]), .IN5(
        N386), .IN6(n786), .Q(n367) );
  AO222X1 U1066 ( .IN1(n784), .IN2(fpTemp[28]), .IN3(n785), .IN4(k[13]), .IN5(
        N387), .IN6(n786), .Q(n366) );
  AO222X1 U1067 ( .IN1(n784), .IN2(fpTemp[29]), .IN3(n785), .IN4(k[14]), .IN5(
        N388), .IN6(n786), .Q(n365) );
  NAND2X0 U1068 ( .IN1(N406), .IN2(n738), .QN(n792) );
  INVX0 U1069 ( .INP(n790), .ZN(n793) );
  NOR4X0 U1070 ( .IN1(n794), .IN2(n795), .IN3(n796), .IN4(n797), .QN(n790) );
  NAND4X0 U1071 ( .IN1(n978), .IN2(n979), .IN3(n980), .IN4(n981), .QN(n797) );
  NAND4X0 U1072 ( .IN1(n982), .IN2(n983), .IN3(n984), .IN4(n989), .QN(n796) );
  NAND3X0 U1073 ( .IN1(n972), .IN2(n973), .IN3(n971), .QN(n795) );
  NAND4X0 U1074 ( .IN1(n974), .IN2(n975), .IN3(n976), .IN4(n977), .QN(n794) );
  NAND2X0 U1075 ( .IN1(n798), .IN2(n799), .QN(n697) );
  AO22X1 U1076 ( .IN1(n800), .IN2(data_in[15]), .IN3(n801), .IN4(
        bestneighborID[15]), .Q(n364) );
  AO22X1 U1077 ( .IN1(n800), .IN2(data_in[14]), .IN3(n801), .IN4(
        bestneighborID[14]), .Q(n363) );
  AO22X1 U1078 ( .IN1(n800), .IN2(data_in[13]), .IN3(n801), .IN4(
        bestneighborID[13]), .Q(n362) );
  AO22X1 U1079 ( .IN1(n800), .IN2(data_in[12]), .IN3(n801), .IN4(
        bestneighborID[12]), .Q(n361) );
  AO221X1 U1080 ( .IN1(n801), .IN2(bestneighborID[11]), .IN3(n802), .IN4(
        data_in[11]), .IN5(n803), .Q(n360) );
  AO221X1 U1081 ( .IN1(n801), .IN2(bestneighborID[10]), .IN3(n802), .IN4(
        data_in[10]), .IN5(n803), .Q(n359) );
  AO221X1 U1082 ( .IN1(n801), .IN2(bestneighborID[9]), .IN3(n802), .IN4(
        data_in[9]), .IN5(n803), .Q(n358) );
  AO221X1 U1083 ( .IN1(n801), .IN2(bestneighborID[8]), .IN3(n802), .IN4(
        data_in[8]), .IN5(n803), .Q(n357) );
  AO221X1 U1084 ( .IN1(n801), .IN2(bestneighborID[7]), .IN3(n802), .IN4(
        data_in[7]), .IN5(n803), .Q(n356) );
  AO221X1 U1085 ( .IN1(n801), .IN2(bestneighborID[6]), .IN3(n802), .IN4(
        data_in[6]), .IN5(n803), .Q(n355) );
  AO221X1 U1086 ( .IN1(n801), .IN2(bestneighborID[5]), .IN3(n802), .IN4(
        data_in[5]), .IN5(n803), .Q(n354) );
  AO221X1 U1087 ( .IN1(n801), .IN2(bestneighborID[4]), .IN3(n802), .IN4(
        data_in[4]), .IN5(n803), .Q(n353) );
  AO221X1 U1088 ( .IN1(n801), .IN2(bestneighborID[3]), .IN3(n802), .IN4(
        data_in[3]), .IN5(n803), .Q(n352) );
  AO221X1 U1089 ( .IN1(n801), .IN2(bestneighborID[2]), .IN3(n802), .IN4(
        data_in[2]), .IN5(n803), .Q(n351) );
  AO221X1 U1090 ( .IN1(n801), .IN2(bestneighborID[1]), .IN3(n802), .IN4(
        data_in[1]), .IN5(n803), .Q(n350) );
  AO22X1 U1091 ( .IN1(n800), .IN2(data_in[0]), .IN3(n801), .IN4(
        bestneighborID[0]), .Q(n349) );
  AO222X1 U1092 ( .IN1(qValue[15]), .IN2(n805), .IN3(n806), .IN4(data_in[15]), 
        .IN5(N456), .IN6(n531), .Q(n348) );
  AO222X1 U1093 ( .IN1(qValue[14]), .IN2(n805), .IN3(n806), .IN4(data_in[14]), 
        .IN5(N455), .IN6(n531), .Q(n347) );
  AO222X1 U1094 ( .IN1(qValue[13]), .IN2(n805), .IN3(n806), .IN4(data_in[13]), 
        .IN5(N454), .IN6(n531), .Q(n346) );
  AO222X1 U1095 ( .IN1(qValue[12]), .IN2(n805), .IN3(n806), .IN4(data_in[12]), 
        .IN5(N453), .IN6(n531), .Q(n345) );
  AO222X1 U1096 ( .IN1(qValue[11]), .IN2(n805), .IN3(n806), .IN4(data_in[11]), 
        .IN5(N452), .IN6(n530), .Q(n344) );
  AO222X1 U1097 ( .IN1(qValue[10]), .IN2(n805), .IN3(n806), .IN4(data_in[10]), 
        .IN5(N451), .IN6(n530), .Q(n343) );
  AO222X1 U1098 ( .IN1(qValue[9]), .IN2(n805), .IN3(n806), .IN4(data_in[9]), 
        .IN5(N450), .IN6(n530), .Q(n342) );
  AO222X1 U1099 ( .IN1(qValue[8]), .IN2(n805), .IN3(n806), .IN4(data_in[8]), 
        .IN5(N449), .IN6(n530), .Q(n341) );
  AO222X1 U1100 ( .IN1(qValue[7]), .IN2(n805), .IN3(n806), .IN4(data_in[7]), 
        .IN5(N448), .IN6(n530), .Q(n340) );
  AO222X1 U1101 ( .IN1(qValue[6]), .IN2(n805), .IN3(n806), .IN4(data_in[6]), 
        .IN5(N447), .IN6(n530), .Q(n339) );
  AO222X1 U1102 ( .IN1(qValue[5]), .IN2(n805), .IN3(n806), .IN4(data_in[5]), 
        .IN5(N446), .IN6(n530), .Q(n338) );
  AO222X1 U1103 ( .IN1(qValue[4]), .IN2(n805), .IN3(n806), .IN4(data_in[4]), 
        .IN5(N445), .IN6(n530), .Q(n337) );
  AO222X1 U1104 ( .IN1(qValue[3]), .IN2(n805), .IN3(n806), .IN4(data_in[3]), 
        .IN5(N444), .IN6(n530), .Q(n336) );
  AO222X1 U1105 ( .IN1(qValue[2]), .IN2(n805), .IN3(n806), .IN4(data_in[2]), 
        .IN5(N443), .IN6(n530), .Q(n335) );
  AO222X1 U1106 ( .IN1(qValue[1]), .IN2(n805), .IN3(n806), .IN4(data_in[1]), 
        .IN5(N442), .IN6(n530), .Q(n334) );
  AO222X1 U1107 ( .IN1(qValue[0]), .IN2(n805), .IN3(n806), .IN4(data_in[0]), 
        .IN5(N441), .IN6(n530), .Q(n333) );
  AO22X1 U1108 ( .IN1(n791), .IN2(done), .IN3(n733), .IN4(nrst), .Q(n332) );
  INVX0 U1109 ( .INP(n722), .ZN(n733) );
  NAND2X0 U1110 ( .IN1(n807), .IN2(n808), .QN(n722) );
  MUX21X1 U1111 ( .IN1(n809), .IN2(wr_en), .S(n810), .Q(n331) );
  AND4X1 U1112 ( .IN1(n696), .IN2(n723), .IN3(n726), .IN4(n811), .Q(n810) );
  NAND2X0 U1113 ( .IN1(n798), .IN2(n808), .QN(n726) );
  NAND2X0 U1114 ( .IN1(n812), .IN2(n807), .QN(n723) );
  OR2X1 U1115 ( .IN1(n800), .IN2(n806), .Q(n809) );
  AO22X1 U1116 ( .IN1(n811), .IN2(betterneighborCount[0]), .IN3(N292), .IN4(
        n814), .Q(n330) );
  AO22X1 U1117 ( .IN1(n811), .IN2(betterneighborCount[1]), .IN3(N293), .IN4(
        n814), .Q(n329) );
  AO22X1 U1118 ( .IN1(n811), .IN2(betterneighborCount[2]), .IN3(N294), .IN4(
        n814), .Q(n328) );
  AO22X1 U1119 ( .IN1(n811), .IN2(betterneighborCount[3]), .IN3(N295), .IN4(
        n814), .Q(n327) );
  AO22X1 U1120 ( .IN1(n811), .IN2(betterneighborCount[4]), .IN3(N296), .IN4(
        n814), .Q(n326) );
  AO22X1 U1121 ( .IN1(n811), .IN2(betterneighborCount[5]), .IN3(N297), .IN4(
        n814), .Q(n325) );
  AO22X1 U1122 ( .IN1(n811), .IN2(betterneighborCount[6]), .IN3(N298), .IN4(
        n814), .Q(n324) );
  AO22X1 U1123 ( .IN1(n811), .IN2(betterneighborCount[7]), .IN3(N299), .IN4(
        n814), .Q(n323) );
  AO22X1 U1124 ( .IN1(n811), .IN2(betterneighborCount[8]), .IN3(N300), .IN4(
        n814), .Q(n322) );
  AO22X1 U1125 ( .IN1(n811), .IN2(betterneighborCount[9]), .IN3(N301), .IN4(
        n814), .Q(n321) );
  AO22X1 U1126 ( .IN1(n811), .IN2(betterneighborCount[10]), .IN3(N302), .IN4(
        n814), .Q(n320) );
  AO22X1 U1127 ( .IN1(n811), .IN2(betterneighborCount[11]), .IN3(N303), .IN4(
        n814), .Q(n319) );
  AO22X1 U1128 ( .IN1(n811), .IN2(betterneighborCount[12]), .IN3(N304), .IN4(
        n814), .Q(n318) );
  AO22X1 U1129 ( .IN1(n811), .IN2(betterneighborCount[13]), .IN3(N305), .IN4(
        n814), .Q(n317) );
  AO22X1 U1130 ( .IN1(n811), .IN2(betterneighborCount[14]), .IN3(N306), .IN4(
        n814), .Q(n316) );
  AO22X1 U1131 ( .IN1(n811), .IN2(betterneighborCount[15]), .IN3(N307), .IN4(
        n814), .Q(n315) );
  AO222X1 U1132 ( .IN1(n816), .IN2(data_out[0]), .IN3(n817), .IN4(N330), .IN5(
        n800), .IN6(betterneighborCount[0]), .Q(n314) );
  AO222X1 U1133 ( .IN1(n816), .IN2(data_out[1]), .IN3(n817), .IN4(N331), .IN5(
        n800), .IN6(betterneighborCount[1]), .Q(n313) );
  AO222X1 U1134 ( .IN1(n816), .IN2(data_out[2]), .IN3(n817), .IN4(i[2]), .IN5(
        n800), .IN6(betterneighborCount[2]), .Q(n312) );
  AO222X1 U1135 ( .IN1(n816), .IN2(data_out[3]), .IN3(n817), .IN4(i[3]), .IN5(
        n800), .IN6(betterneighborCount[3]), .Q(n311) );
  AO222X1 U1136 ( .IN1(n816), .IN2(data_out[4]), .IN3(n817), .IN4(i[4]), .IN5(
        n800), .IN6(betterneighborCount[4]), .Q(n310) );
  AO222X1 U1137 ( .IN1(n816), .IN2(data_out[5]), .IN3(n817), .IN4(i[5]), .IN5(
        n800), .IN6(betterneighborCount[5]), .Q(n309) );
  AO222X1 U1138 ( .IN1(n816), .IN2(data_out[6]), .IN3(n817), .IN4(i[6]), .IN5(
        n800), .IN6(betterneighborCount[6]), .Q(n308) );
  AO222X1 U1139 ( .IN1(n816), .IN2(data_out[7]), .IN3(n817), .IN4(i[7]), .IN5(
        n800), .IN6(betterneighborCount[7]), .Q(n307) );
  AO222X1 U1140 ( .IN1(n816), .IN2(data_out[8]), .IN3(n817), .IN4(i[8]), .IN5(
        n800), .IN6(betterneighborCount[8]), .Q(n306) );
  AO222X1 U1141 ( .IN1(n816), .IN2(data_out[9]), .IN3(n817), .IN4(i[9]), .IN5(
        n800), .IN6(betterneighborCount[9]), .Q(n305) );
  AO222X1 U1142 ( .IN1(n816), .IN2(data_out[10]), .IN3(n817), .IN4(i[10]), 
        .IN5(n800), .IN6(betterneighborCount[10]), .Q(n304) );
  AO222X1 U1143 ( .IN1(n816), .IN2(data_out[11]), .IN3(n817), .IN4(i[11]), 
        .IN5(n800), .IN6(betterneighborCount[11]), .Q(n303) );
  AO222X1 U1144 ( .IN1(n816), .IN2(data_out[12]), .IN3(n817), .IN4(i[12]), 
        .IN5(n800), .IN6(betterneighborCount[12]), .Q(n302) );
  AO222X1 U1145 ( .IN1(n816), .IN2(data_out[13]), .IN3(n817), .IN4(i[13]), 
        .IN5(n800), .IN6(betterneighborCount[13]), .Q(n301) );
  AO222X1 U1146 ( .IN1(n816), .IN2(data_out[14]), .IN3(n817), .IN4(i[14]), 
        .IN5(n800), .IN6(betterneighborCount[14]), .Q(n300) );
  AO222X1 U1147 ( .IN1(n816), .IN2(data_out[15]), .IN3(n817), .IN4(i[15]), 
        .IN5(n800), .IN6(betterneighborCount[15]), .Q(n299) );
  NAND2X0 U1148 ( .IN1(n818), .IN2(nrst), .QN(n813) );
  NAND3X0 U1149 ( .IN1(n696), .IN2(n819), .IN3(nrst), .QN(n718) );
  AO22X1 U1150 ( .IN1(n820), .IN2(bestvalue[0]), .IN3(n821), .IN4(N441), .Q(
        n298) );
  NAND2X0 U1151 ( .IN1(n822), .IN2(n823), .QN(n297) );
  MUX21X1 U1152 ( .IN1(n970), .IN2(n986), .S(n824), .Q(n822) );
  AO22X1 U1153 ( .IN1(n820), .IN2(N164), .IN3(n821), .IN4(N331), .Q(n296) );
  AO22X1 U1154 ( .IN1(n820), .IN2(besthop[2]), .IN3(n821), .IN4(i[2]), .Q(n295) );
  AO22X1 U1155 ( .IN1(n820), .IN2(besthop[3]), .IN3(n821), .IN4(i[3]), .Q(n294) );
  AO22X1 U1156 ( .IN1(n820), .IN2(besthop[4]), .IN3(n821), .IN4(i[4]), .Q(n293) );
  AO22X1 U1157 ( .IN1(n820), .IN2(besthop[5]), .IN3(n821), .IN4(i[5]), .Q(n292) );
  NAND2X0 U1158 ( .IN1(n825), .IN2(n823), .QN(n291) );
  MUX21X1 U1159 ( .IN1(n969), .IN2(n985), .S(n824), .Q(n825) );
  AO22X1 U1160 ( .IN1(n820), .IN2(besthop[7]), .IN3(n821), .IN4(i[7]), .Q(n290) );
  AO22X1 U1161 ( .IN1(n820), .IN2(besthop[8]), .IN3(n821), .IN4(i[8]), .Q(n289) );
  AO22X1 U1162 ( .IN1(n820), .IN2(besthop[9]), .IN3(n821), .IN4(i[9]), .Q(n288) );
  NOR2X0 U1163 ( .IN1(n990), .IN2(n826), .QN(n287) );
  AO22X1 U1164 ( .IN1(n827), .IN2(address[1]), .IN3(nrst), .IN4(n828), .Q(n286) );
  OR4X1 U1165 ( .IN1(n829), .IN2(n830), .IN3(n831), .IN4(n832), .Q(n828) );
  AO222X1 U1166 ( .IN1(N501), .IN2(n754), .IN3(N319), .IN4(n815), .IN5(N163), 
        .IN6(n833), .Q(n832) );
  AO221X1 U1167 ( .IN1(N150), .IN2(n834), .IN3(N330), .IN4(n835), .IN5(n751), 
        .Q(n831) );
  INVX0 U1168 ( .INP(n708), .ZN(n751) );
  AO222X1 U1169 ( .IN1(N472), .IN2(n746), .IN3(N150), .IN4(n836), .IN5(N418), 
        .IN6(n738), .Q(n830) );
  AO222X1 U1170 ( .IN1(N330), .IN2(n837), .IN3(N330), .IN4(n737), .IN5(N150), 
        .IN6(n838), .Q(n829) );
  AO22X1 U1171 ( .IN1(n827), .IN2(address[2]), .IN3(nrst), .IN4(n839), .Q(n285) );
  OR4X1 U1172 ( .IN1(n840), .IN2(n841), .IN3(n842), .IN4(n843), .Q(n839) );
  AO222X1 U1173 ( .IN1(N502), .IN2(n754), .IN3(N320), .IN4(n815), .IN5(N164), 
        .IN6(n833), .Q(n843) );
  AO221X1 U1174 ( .IN1(N151), .IN2(n834), .IN3(N331), .IN4(n835), .IN5(n802), 
        .Q(n842) );
  AO222X1 U1175 ( .IN1(N473), .IN2(n746), .IN3(N151), .IN4(n836), .IN5(N419), 
        .IN6(n738), .Q(n841) );
  AO222X1 U1176 ( .IN1(N331), .IN2(n837), .IN3(N331), .IN4(n737), .IN5(N151), 
        .IN6(n838), .Q(n840) );
  MUX21X1 U1177 ( .IN1(address[3]), .IN2(n844), .S(n826), .Q(n284) );
  OR4X1 U1178 ( .IN1(n845), .IN2(n846), .IN3(n847), .IN4(n848), .Q(n844) );
  AO222X1 U1179 ( .IN1(N165), .IN2(n833), .IN3(N503), .IN4(n754), .IN5(N332), 
        .IN6(n737), .Q(n848) );
  AO221X1 U1180 ( .IN1(N332), .IN2(n835), .IN3(N321), .IN4(n815), .IN5(n849), 
        .Q(n847) );
  AO21X1 U1181 ( .IN1(N230), .IN2(n834), .IN3(n748), .Q(n849) );
  AO221X1 U1182 ( .IN1(N474), .IN2(n746), .IN3(N420), .IN4(n738), .IN5(n730), 
        .Q(n846) );
  AO222X1 U1183 ( .IN1(N230), .IN2(n838), .IN3(N332), .IN4(n837), .IN5(N230), 
        .IN6(n836), .Q(n845) );
  AO22X1 U1184 ( .IN1(n827), .IN2(address[4]), .IN3(nrst), .IN4(n850), .Q(n283) );
  OR4X1 U1185 ( .IN1(n851), .IN2(n852), .IN3(n853), .IN4(n854), .Q(n850) );
  AO222X1 U1186 ( .IN1(N166), .IN2(n833), .IN3(N504), .IN4(n754), .IN5(N188), 
        .IN6(n737), .Q(n854) );
  AO222X1 U1187 ( .IN1(N267), .IN2(n835), .IN3(N153), .IN4(n834), .IN5(N322), 
        .IN6(n815), .Q(n853) );
  AO22X1 U1188 ( .IN1(N421), .IN2(n738), .IN3(N475), .IN4(n746), .Q(n852) );
  AO222X1 U1189 ( .IN1(N534), .IN2(n838), .IN3(N333), .IN4(n837), .IN5(N231), 
        .IN6(n836), .Q(n851) );
  AO22X1 U1190 ( .IN1(n827), .IN2(address[5]), .IN3(nrst), .IN4(n855), .Q(n282) );
  OR4X1 U1191 ( .IN1(n856), .IN2(n857), .IN3(n858), .IN4(n859), .Q(n855) );
  AO222X1 U1192 ( .IN1(N167), .IN2(n833), .IN3(N505), .IN4(n754), .IN5(N189), 
        .IN6(n737), .Q(n859) );
  AO222X1 U1193 ( .IN1(N268), .IN2(n835), .IN3(N154), .IN4(n834), .IN5(N323), 
        .IN6(n815), .Q(n858) );
  AO22X1 U1194 ( .IN1(N422), .IN2(n738), .IN3(N476), .IN4(n746), .Q(n857) );
  AO222X1 U1195 ( .IN1(N535), .IN2(n838), .IN3(N334), .IN4(n837), .IN5(N232), 
        .IN6(n836), .Q(n856) );
  AO22X1 U1196 ( .IN1(n827), .IN2(address[6]), .IN3(nrst), .IN4(n860), .Q(n281) );
  OR4X1 U1197 ( .IN1(n861), .IN2(n862), .IN3(n863), .IN4(n864), .Q(n860) );
  AO222X1 U1198 ( .IN1(N506), .IN2(n754), .IN3(N324), .IN4(n815), .IN5(N168), 
        .IN6(n833), .Q(n864) );
  AO221X1 U1199 ( .IN1(N155), .IN2(n834), .IN3(N269), .IN4(n835), .IN5(n748), 
        .Q(n863) );
  AO222X1 U1200 ( .IN1(N477), .IN2(n746), .IN3(N233), .IN4(n836), .IN5(N423), 
        .IN6(n738), .Q(n862) );
  AO222X1 U1201 ( .IN1(N335), .IN2(n837), .IN3(N190), .IN4(n737), .IN5(N536), 
        .IN6(n838), .Q(n861) );
  MUX21X1 U1202 ( .IN1(address[7]), .IN2(n865), .S(n826), .Q(n280) );
  OR4X1 U1203 ( .IN1(n866), .IN2(n867), .IN3(n868), .IN4(n869), .Q(n865) );
  AO222X1 U1204 ( .IN1(N169), .IN2(n833), .IN3(N507), .IN4(n754), .IN5(N191), 
        .IN6(n737), .Q(n869) );
  AO221X1 U1205 ( .IN1(N270), .IN2(n835), .IN3(N325), .IN4(n815), .IN5(n870), 
        .Q(n868) );
  AO21X1 U1206 ( .IN1(N156), .IN2(n834), .IN3(n748), .Q(n870) );
  INVX0 U1207 ( .INP(n747), .ZN(n748) );
  AO221X1 U1208 ( .IN1(N478), .IN2(n746), .IN3(N424), .IN4(n738), .IN5(n730), 
        .Q(n867) );
  AO222X1 U1209 ( .IN1(N537), .IN2(n838), .IN3(N336), .IN4(n837), .IN5(N234), 
        .IN6(n836), .Q(n866) );
  AO22X1 U1210 ( .IN1(n827), .IN2(address[8]), .IN3(nrst), .IN4(n871), .Q(n279) );
  OR4X1 U1211 ( .IN1(n872), .IN2(n873), .IN3(n874), .IN4(n875), .Q(n871) );
  AO222X1 U1212 ( .IN1(N170), .IN2(n833), .IN3(N508), .IN4(n754), .IN5(N192), 
        .IN6(n737), .Q(n875) );
  AO222X1 U1213 ( .IN1(N271), .IN2(n835), .IN3(N157), .IN4(n834), .IN5(N326), 
        .IN6(n815), .Q(n874) );
  AO22X1 U1214 ( .IN1(N425), .IN2(n738), .IN3(N479), .IN4(n746), .Q(n873) );
  AO222X1 U1215 ( .IN1(N538), .IN2(n838), .IN3(N337), .IN4(n837), .IN5(N235), 
        .IN6(n836), .Q(n872) );
  INVX0 U1216 ( .INP(n826), .ZN(n827) );
  MUX21X1 U1217 ( .IN1(address[9]), .IN2(n876), .S(n826), .Q(n278) );
  OR4X1 U1218 ( .IN1(n877), .IN2(n878), .IN3(n879), .IN4(n880), .Q(n876) );
  AO222X1 U1219 ( .IN1(N171), .IN2(n833), .IN3(N509), .IN4(n754), .IN5(N193), 
        .IN6(n737), .Q(n880) );
  AO222X1 U1220 ( .IN1(N272), .IN2(n835), .IN3(N158), .IN4(n834), .IN5(N327), 
        .IN6(n815), .Q(n879) );
  AO221X1 U1221 ( .IN1(N480), .IN2(n746), .IN3(N426), .IN4(n738), .IN5(n730), 
        .Q(n878) );
  AO222X1 U1222 ( .IN1(N539), .IN2(n838), .IN3(N338), .IN4(n837), .IN5(N236), 
        .IN6(n836), .Q(n877) );
  MUX21X1 U1223 ( .IN1(address[10]), .IN2(n881), .S(n826), .Q(n277) );
  NAND4X0 U1224 ( .IN1(n805), .IN2(n882), .IN3(n758), .IN4(n883), .QN(n826) );
  AND3X1 U1225 ( .IN1(n745), .IN2(n747), .IN3(n708), .Q(n883) );
  NAND2X0 U1226 ( .IN1(n808), .IN2(n884), .QN(n747) );
  NOR3X0 U1227 ( .IN1(n885), .IN2(n707), .IN3(n755), .QN(n758) );
  INVX0 U1228 ( .INP(n706), .ZN(n882) );
  NAND3X0 U1229 ( .IN1(n696), .IN2(n695), .IN3(n886), .QN(n706) );
  NAND3X0 U1230 ( .IN1(n887), .IN2(n884), .IN3(start), .QN(n886) );
  OR4X1 U1231 ( .IN1(n888), .IN2(n889), .IN3(n890), .IN4(n891), .Q(n881) );
  AO222X1 U1232 ( .IN1(N172), .IN2(n833), .IN3(N510), .IN4(n754), .IN5(N194), 
        .IN6(n737), .Q(n891) );
  AND2X1 U1233 ( .IN1(N160), .IN2(n759), .Q(n833) );
  NAND3X0 U1234 ( .IN1(n700), .IN2(n727), .IN3(n698), .QN(n759) );
  INVX0 U1235 ( .INP(n892), .ZN(n700) );
  AO222X1 U1236 ( .IN1(N273), .IN2(n835), .IN3(N159), .IN4(n834), .IN5(N328), 
        .IN6(n815), .Q(n890) );
  NAND2X0 U1237 ( .IN1(n818), .IN2(n893), .QN(n819) );
  INVX0 U1238 ( .INP(n735), .ZN(n818) );
  NAND2X0 U1239 ( .IN1(N130), .IN2(n885), .QN(n698) );
  INVX0 U1240 ( .INP(n725), .ZN(n885) );
  NAND2X0 U1241 ( .IN1(n799), .IN2(n884), .QN(n725) );
  NAND2X0 U1242 ( .IN1(n707), .IN2(n894), .QN(n702) );
  INVX0 U1243 ( .INP(n724), .ZN(n707) );
  AO221X1 U1244 ( .IN1(N481), .IN2(n746), .IN3(N427), .IN4(n738), .IN5(n730), 
        .Q(n889) );
  NAND4X0 U1245 ( .IN1(n804), .IN2(n895), .IN3(n708), .IN4(n696), .QN(n730) );
  NAND2X0 U1246 ( .IN1(n887), .IN2(n807), .QN(n696) );
  NAND2X0 U1247 ( .IN1(n812), .IN2(n884), .QN(n708) );
  NAND2X0 U1248 ( .IN1(n887), .IN2(n884), .QN(n895) );
  NOR2X0 U1249 ( .IN1(state[3]), .IN2(state[2]), .QN(n884) );
  INVX0 U1250 ( .INP(n762), .ZN(n804) );
  NAND2X0 U1251 ( .IN1(n896), .IN2(n887), .QN(n695) );
  NAND2X0 U1252 ( .IN1(n896), .IN2(n808), .QN(n745) );
  NOR2X0 U1253 ( .IN1(n897), .IN2(state[0]), .QN(n808) );
  AO222X1 U1254 ( .IN1(N540), .IN2(n838), .IN3(N339), .IN4(n837), .IN5(N237), 
        .IN6(n836), .Q(n888) );
  NAND2X0 U1255 ( .IN1(n892), .IN2(n699), .QN(n709) );
  INVX0 U1256 ( .INP(N160), .ZN(n699) );
  NOR2X0 U1257 ( .IN1(n894), .IN2(n724), .QN(n892) );
  NAND2X0 U1258 ( .IN1(n798), .IN2(n887), .QN(n724) );
  NOR2X0 U1259 ( .IN1(state[1]), .IN2(state[0]), .QN(n887) );
  NAND4X0 U1260 ( .IN1(n898), .IN2(n899), .IN3(n900), .IN4(n901), .QN(n894) );
  NOR4X0 U1261 ( .IN1(data_in[9]), .IN2(data_in[15]), .IN3(data_in[14]), .IN4(
        data_in[13]), .QN(n901) );
  OA21X1 U1262 ( .IN1(n902), .IN2(n903), .IN3(n904), .Q(n900) );
  OA21X1 U1263 ( .IN1(n905), .IN2(n906), .IN3(n907), .Q(n902) );
  AND3X1 U1264 ( .IN1(n908), .IN2(n909), .IN3(n910), .Q(n905) );
  OA21X1 U1265 ( .IN1(n735), .IN2(n893), .IN3(n736), .Q(n691) );
  AO21X1 U1266 ( .IN1(mybest[15]), .IN2(n911), .IN3(n912), .Q(n893) );
  OA22X1 U1267 ( .IN1(mybest[15]), .IN2(n911), .IN3(n913), .IN4(n914), .Q(n912) );
  AND2X1 U1268 ( .IN1(n915), .IN2(mybest[14]), .Q(n914) );
  OA221X1 U1269 ( .IN1(mybest[13]), .IN2(n916), .IN3(mybest[14]), .IN4(n915), 
        .IN5(n917), .Q(n913) );
  AO221X1 U1270 ( .IN1(mybest[12]), .IN2(n899), .IN3(mybest[13]), .IN4(n916), 
        .IN5(n918), .Q(n917) );
  OA221X1 U1271 ( .IN1(mybest[11]), .IN2(n898), .IN3(mybest[12]), .IN4(n899), 
        .IN5(n919), .Q(n918) );
  AO221X1 U1272 ( .IN1(mybest[10]), .IN2(n904), .IN3(mybest[11]), .IN4(n898), 
        .IN5(n920), .Q(n919) );
  OA221X1 U1273 ( .IN1(mybest[9]), .IN2(n921), .IN3(mybest[10]), .IN4(n904), 
        .IN5(n922), .Q(n920) );
  AO221X1 U1274 ( .IN1(mybest[8]), .IN2(n903), .IN3(mybest[9]), .IN4(n921), 
        .IN5(n923), .Q(n922) );
  OA221X1 U1275 ( .IN1(mybest[7]), .IN2(n907), .IN3(mybest[8]), .IN4(n903), 
        .IN5(n924), .Q(n923) );
  AO221X1 U1276 ( .IN1(mybest[6]), .IN2(n906), .IN3(mybest[7]), .IN4(n907), 
        .IN5(n925), .Q(n924) );
  OA221X1 U1277 ( .IN1(mybest[5]), .IN2(n909), .IN3(mybest[6]), .IN4(n906), 
        .IN5(n926), .Q(n925) );
  AO221X1 U1278 ( .IN1(mybest[4]), .IN2(n910), .IN3(mybest[5]), .IN4(n909), 
        .IN5(n927), .Q(n926) );
  OA221X1 U1279 ( .IN1(mybest[3]), .IN2(n908), .IN3(mybest[4]), .IN4(n910), 
        .IN5(n928), .Q(n927) );
  AO222X1 U1280 ( .IN1(n929), .IN2(n930), .IN3(mybest[2]), .IN4(n931), .IN5(
        mybest[3]), .IN6(n908), .Q(n928) );
  OR2X1 U1281 ( .IN1(n930), .IN2(n929), .Q(n931) );
  INVX0 U1282 ( .INP(data_in[2]), .ZN(n930) );
  OA22X1 U1283 ( .IN1(mybest[1]), .IN2(n932), .IN3(n933), .IN4(n934), .Q(n929)
         );
  AO21X1 U1284 ( .IN1(mybest[1]), .IN2(n932), .IN3(mybest[0]), .Q(n934) );
  INVX0 U1285 ( .INP(data_in[0]), .ZN(n933) );
  INVX0 U1286 ( .INP(data_in[1]), .ZN(n932) );
  INVX0 U1287 ( .INP(data_in[3]), .ZN(n908) );
  INVX0 U1288 ( .INP(data_in[4]), .ZN(n910) );
  INVX0 U1289 ( .INP(data_in[5]), .ZN(n909) );
  INVX0 U1290 ( .INP(data_in[6]), .ZN(n906) );
  INVX0 U1291 ( .INP(data_in[7]), .ZN(n907) );
  INVX0 U1292 ( .INP(data_in[8]), .ZN(n903) );
  INVX0 U1293 ( .INP(data_in[9]), .ZN(n921) );
  INVX0 U1294 ( .INP(data_in[10]), .ZN(n904) );
  INVX0 U1295 ( .INP(data_in[11]), .ZN(n898) );
  INVX0 U1296 ( .INP(data_in[12]), .ZN(n899) );
  INVX0 U1297 ( .INP(data_in[14]), .ZN(n915) );
  INVX0 U1298 ( .INP(data_in[13]), .ZN(n916) );
  INVX0 U1299 ( .INP(data_in[15]), .ZN(n911) );
  NAND2X0 U1300 ( .IN1(n812), .IN2(n798), .QN(n735) );
  NOR2X0 U1301 ( .IN1(n935), .IN2(state[3]), .QN(n798) );
  NAND2X0 U1302 ( .IN1(N511), .IN2(n755), .QN(n727) );
  INVX0 U1303 ( .INP(n714), .ZN(n755) );
  NAND2X0 U1304 ( .IN1(n896), .IN2(n799), .QN(n714) );
  AO22X1 U1305 ( .IN1(n820), .IN2(besthop[10]), .IN3(n821), .IN4(i[10]), .Q(
        n276) );
  AO22X1 U1306 ( .IN1(n820), .IN2(besthop[11]), .IN3(n821), .IN4(i[11]), .Q(
        n275) );
  AO22X1 U1307 ( .IN1(n820), .IN2(besthop[12]), .IN3(n821), .IN4(i[12]), .Q(
        n274) );
  AO22X1 U1308 ( .IN1(n820), .IN2(besthop[13]), .IN3(n821), .IN4(i[13]), .Q(
        n273) );
  AO22X1 U1309 ( .IN1(n820), .IN2(besthop[14]), .IN3(n821), .IN4(i[14]), .Q(
        n272) );
  AO22X1 U1310 ( .IN1(n820), .IN2(besthop[15]), .IN3(n821), .IN4(i[15]), .Q(
        n271) );
  NAND2X0 U1311 ( .IN1(n936), .IN2(n823), .QN(n270) );
  MUX21X1 U1312 ( .IN1(n968), .IN2(n649), .S(n824), .Q(n936) );
  NAND2X0 U1313 ( .IN1(n937), .IN2(n823), .QN(n269) );
  MUX21X1 U1314 ( .IN1(n967), .IN2(n650), .S(n824), .Q(n937) );
  NAND2X0 U1315 ( .IN1(n938), .IN2(n823), .QN(n268) );
  MUX21X1 U1316 ( .IN1(n966), .IN2(n651), .S(n824), .Q(n938) );
  NAND2X0 U1317 ( .IN1(n939), .IN2(n823), .QN(n267) );
  MUX21X1 U1318 ( .IN1(n965), .IN2(n652), .S(n824), .Q(n939) );
  NAND2X0 U1319 ( .IN1(n940), .IN2(n823), .QN(n266) );
  MUX21X1 U1320 ( .IN1(n653), .IN2(n964), .S(n820), .Q(n940) );
  NAND2X0 U1321 ( .IN1(n941), .IN2(n823), .QN(n265) );
  MUX21X1 U1322 ( .IN1(n654), .IN2(n963), .S(n820), .Q(n941) );
  NAND2X0 U1323 ( .IN1(n942), .IN2(n823), .QN(n264) );
  MUX21X1 U1324 ( .IN1(n655), .IN2(n962), .S(n820), .Q(n942) );
  NAND2X0 U1325 ( .IN1(n943), .IN2(n823), .QN(n263) );
  MUX21X1 U1326 ( .IN1(n961), .IN2(n656), .S(n824), .Q(n943) );
  NAND2X0 U1327 ( .IN1(n944), .IN2(n823), .QN(n262) );
  MUX21X1 U1328 ( .IN1(n960), .IN2(n657), .S(n824), .Q(n944) );
  NAND2X0 U1329 ( .IN1(n945), .IN2(n823), .QN(n261) );
  MUX21X1 U1330 ( .IN1(n959), .IN2(n658), .S(n824), .Q(n945) );
  NAND2X0 U1331 ( .IN1(n946), .IN2(n823), .QN(n260) );
  MUX21X1 U1332 ( .IN1(n958), .IN2(n659), .S(n824), .Q(n946) );
  NAND2X0 U1333 ( .IN1(n947), .IN2(n823), .QN(n259) );
  MUX21X1 U1334 ( .IN1(n957), .IN2(n660), .S(n824), .Q(n947) );
  NAND2X0 U1335 ( .IN1(n948), .IN2(n823), .QN(n258) );
  MUX21X1 U1336 ( .IN1(n956), .IN2(n661), .S(n824), .Q(n948) );
  NAND2X0 U1337 ( .IN1(n949), .IN2(n823), .QN(n257) );
  MUX21X1 U1338 ( .IN1(n955), .IN2(n662), .S(n824), .Q(n949) );
  NAND2X0 U1339 ( .IN1(n950), .IN2(n823), .QN(n256) );
  MUX21X1 U1340 ( .IN1(n954), .IN2(n663), .S(n824), .Q(n950) );
  NAND2X0 U1341 ( .IN1(n736), .IN2(n791), .QN(n783) );
  INVX0 U1342 ( .INP(n742), .ZN(n791) );
  NAND2X0 U1343 ( .IN1(n812), .IN2(n896), .QN(n736) );
  NOR2X0 U1344 ( .IN1(n951), .IN2(state[2]), .QN(n896) );
  NOR2X0 U1345 ( .IN1(n952), .IN2(state[1]), .QN(n812) );
  OA21X1 U1346 ( .IN1(n741), .IN2(en), .IN3(n762), .Q(n742) );
  NAND2X0 U1347 ( .IN1(nrst), .IN2(n715), .QN(n762) );
  NAND2X0 U1348 ( .IN1(n807), .IN2(n799), .QN(n715) );
  NOR2X0 U1349 ( .IN1(n952), .IN2(n897), .QN(n799) );
  NOR2X0 U1350 ( .IN1(n951), .IN2(n935), .QN(n807) );
  NAND2X0 U1351 ( .IN1(n987), .IN2(n953), .QN(N419) );
  NAND2X0 U1352 ( .IN1(n988), .IN2(n953), .QN(N413) );
  INVX0 U1353 ( .INP(N406), .ZN(n953) );
  NOR2X0 U1354 ( .IN1(n62), .IN2(N406), .QN(N418) );
  NOR2X0 U1355 ( .IN1(n61), .IN2(N406), .QN(N1276) );
  NOR2X0 U1356 ( .IN1(n60), .IN2(N406), .QN(N1272) );
  NOR2X0 U1357 ( .IN1(n59), .IN2(N406), .QN(N1270) );
  NOR2X0 U1358 ( .IN1(n58), .IN2(N406), .QN(N1268) );
  NOR2X0 U1359 ( .IN1(n57), .IN2(N406), .QN(N1266) );
  NOR2X0 U1360 ( .IN1(n56), .IN2(N406), .QN(N1264) );
  NOR2X0 U1361 ( .IN1(n55), .IN2(N406), .QN(N1262) );
endmodule

