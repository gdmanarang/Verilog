
module fixSinkList_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_2 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_3 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_inc_4 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module fixSinkList_DW01_add_11 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [15:1] carry;

  FADDX1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .S(SUM[15]) );
  FADDX1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FADDX1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FADDX1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FADDX1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FADDX1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FADDX1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FADDX1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8])
         );
  FADDX1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7])
         );
  FADDX1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6])
         );
  FADDX1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5])
         );
  FADDX1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4])
         );
  FADDX1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3])
         );
  FADDX1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2])
         );
  FADDX1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n1), .CO(carry[2]), .S(SUM[1]) );
  AND2X1 U1 ( .IN1(B[0]), .IN2(A[0]), .Q(n1) );
  XOR2X1 U2 ( .IN1(B[0]), .IN2(A[0]), .Q(SUM[0]) );
endmodule


module fixSinkList ( clock, nrst, en, start, address, wr_en, data_in, data_out, 
        done );
  output [10:0] address;
  input [15:0] data_in;
  output [15:0] data_out;
  input clock, nrst, en, start;
  output wr_en, done;
  wire   N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N119,
         N120, N121, N122, N123, N124, N125, N126, N127, N128, N133, N134,
         N135, N136, N137, N138, N139, N141, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N152, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N193, N194, N195, N196, N197, N198, N199,
         N200, N201, N202, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N259, N260, N261, N262, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N357, N358, N359, N360, N361, N362,
         N363, N368, N369, N370, N371, N372, N373, N374, N391, N392, N393,
         N394, N395, N396, N397, N398, N399, N400, N401, N402, N403, N404,
         N405, N406, N407, N408, N409, N410, N411, N412, N413, N414, N415,
         N416, N417, N418, N419, N420, N421, N422, N476, N477, N478, N479,
         N480, N481, N482, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, n71, n79, n80, n81, n84, n89, n90, n91, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, N390, N389, N388, N387, N386, N385,
         N384, N383, N382, N381, N380, N379, N378, N377, N376, N375,
         \add_160/carry[10] , \add_160/carry[9] , \add_160/carry[8] ,
         \add_160/carry[7] , \add_160/carry[6] , \add_160/carry[5] ,
         \add_160/carry[4] , \add_160/carry[3] , \add_155/carry[10] ,
         \add_155/carry[9] , \add_155/carry[8] , \add_155/carry[7] ,
         \add_155/carry[6] , \add_155/carry[5] , \add_121/carry[10] ,
         \add_121/carry[9] , \add_121/carry[8] , \add_121/carry[7] ,
         \add_121/carry[6] , \add_121/carry[5] , \add_115/carry[10] ,
         \add_115/carry[9] , \add_115/carry[8] , \add_115/carry[7] ,
         \add_115/carry[6] , \add_115/carry[5] , \add_92/carry[10] ,
         \add_92/carry[9] , \add_92/carry[8] , \add_92/carry[7] ,
         \add_92/carry[6] , \add_92/carry[5] , \add_92/carry[4] ,
         \add_92/carry[3] , \add_87/carry[10] , \add_87/carry[9] ,
         \add_87/carry[8] , \add_87/carry[7] , \add_87/carry[6] ,
         \add_87/carry[5] , \add_0_root_add_67_2/carry[10] ,
         \add_0_root_add_67_2/carry[9] , \add_0_root_add_67_2/carry[8] ,
         \add_0_root_add_67_2/carry[7] , \add_0_root_add_67_2/carry[6] ,
         \add_0_root_add_67_2/carry[5] , \add_55/carry[10] , \add_55/carry[9] ,
         \add_55/carry[8] , \add_55/carry[7] , \add_55/carry[6] ,
         \add_55/carry[5] , \r241/carry[10] , \r241/carry[9] , \r241/carry[8] ,
         \r241/carry[7] , \r241/carry[6] , \r241/carry[5] , \r230/carry[10] ,
         \r230/carry[9] , \r230/carry[8] , \r229/carry[10] , \r229/carry[9] ,
         \r229/carry[8] , \r229/carry[7] , \r229/carry[6] , \r229/carry[5] ,
         \r229/carry[4] , \r229/carry[3] , n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510;
  wire   [3:0] state;
  wire   [15:0] j;
  wire   [15:0] i;
  wire   [15:0] k;
  wire   [15:0] knownSinkCount;
  wire   [15:0] neighborCount;
  wire   [15:0] knownSinks;
  wire   [15:0] sinkIDCount;
  wire   [15:0] worstHops;

  DFFX1 \state_reg[1]  ( .D(n388), .CLK(clock), .Q(state[1]), .QN(n80) );
  DFFX1 \state_reg[2]  ( .D(n387), .CLK(clock), .Q(state[2]), .QN(n79) );
  DFFX1 \state_reg[3]  ( .D(n389), .CLK(clock), .Q(state[3]), .QN(n71) );
  DFFSSRX1 \state_reg[0]  ( .D(nrst), .RSTB(n217), .SETB(n495), .CLK(clock), 
        .Q(state[0]), .QN(n81) );
  AO22X1 U80 ( .IN1(n96), .IN2(n97), .IN3(address[1]), .IN4(n493), .Q(n232) );
  OR4X1 U81 ( .IN1(n98), .IN2(n99), .IN3(n100), .IN4(n101), .Q(n96) );
  AO222X1 U82 ( .IN1(N193), .IN2(n90), .IN3(N193), .IN4(n95), .IN5(N309), 
        .IN6(n91), .Q(n101) );
  AO221X1 U83 ( .IN1(N205), .IN2(n94), .IN3(N205), .IN4(n93), .IN5(n102), .Q(
        n100) );
  AO221X1 U84 ( .IN1(N141), .IN2(n503), .IN3(N108), .IN4(n501), .IN5(n492), 
        .Q(n99) );
  AO222X1 U85 ( .IN1(N133), .IN2(n509), .IN3(N119), .IN4(n89), .IN5(N108), 
        .IN6(n507), .Q(n98) );
  AO22X1 U86 ( .IN1(address[2]), .IN2(n493), .IN3(n84), .IN4(n105), .Q(n233)
         );
  OR2X1 U87 ( .IN1(n106), .IN2(n107), .Q(n105) );
  AO221X1 U88 ( .IN1(N142), .IN2(n503), .IN3(N109), .IN4(n501), .IN5(n108), 
        .Q(n107) );
  AO222X1 U89 ( .IN1(N134), .IN2(n509), .IN3(N120), .IN4(n89), .IN5(N109), 
        .IN6(n507), .Q(n108) );
  AO221X1 U90 ( .IN1(N194), .IN2(n90), .IN3(N310), .IN4(n91), .IN5(n109), .Q(
        n106) );
  AO222X1 U91 ( .IN1(N486), .IN2(n93), .IN3(N206), .IN4(n94), .IN5(N194), 
        .IN6(n95), .Q(n109) );
  AO22X1 U92 ( .IN1(n110), .IN2(n97), .IN3(address[3]), .IN4(n493), .Q(n234)
         );
  OR4X1 U93 ( .IN1(n111), .IN2(n112), .IN3(n113), .IN4(n114), .Q(n110) );
  AO222X1 U94 ( .IN1(N311), .IN2(n91), .IN3(N195), .IN4(n90), .IN5(N121), 
        .IN6(n89), .Q(n114) );
  AO222X1 U95 ( .IN1(N487), .IN2(n93), .IN3(N207), .IN4(n94), .IN5(N195), 
        .IN6(n95), .Q(n113) );
  AO21X1 U96 ( .IN1(N110), .IN2(n501), .IN3(n115), .Q(n112) );
  AO222X1 U97 ( .IN1(N110), .IN2(n507), .IN3(N135), .IN4(n509), .IN5(N143), 
        .IN6(n503), .Q(n111) );
  AO22X1 U98 ( .IN1(address[4]), .IN2(n493), .IN3(n84), .IN4(n116), .Q(n235)
         );
  OR2X1 U99 ( .IN1(n117), .IN2(n118), .Q(n116) );
  AO221X1 U100 ( .IN1(N144), .IN2(n503), .IN3(N111), .IN4(n501), .IN5(n119), 
        .Q(n118) );
  AO222X1 U101 ( .IN1(N368), .IN2(n509), .IN3(N122), .IN4(n89), .IN5(N357), 
        .IN6(n507), .Q(n119) );
  AO221X1 U102 ( .IN1(N476), .IN2(n90), .IN3(N312), .IN4(n91), .IN5(n120), .Q(
        n117) );
  AO222X1 U103 ( .IN1(N488), .IN2(n93), .IN3(N208), .IN4(n94), .IN5(N196), 
        .IN6(n95), .Q(n120) );
  AO22X1 U104 ( .IN1(address[5]), .IN2(n493), .IN3(n84), .IN4(n121), .Q(n236)
         );
  OR2X1 U105 ( .IN1(n122), .IN2(n123), .Q(n121) );
  AO221X1 U106 ( .IN1(N145), .IN2(n503), .IN3(N112), .IN4(n501), .IN5(n124), 
        .Q(n123) );
  AO222X1 U107 ( .IN1(N369), .IN2(n509), .IN3(N123), .IN4(n89), .IN5(N358), 
        .IN6(n507), .Q(n124) );
  AO221X1 U108 ( .IN1(N477), .IN2(n90), .IN3(N313), .IN4(n91), .IN5(n125), .Q(
        n122) );
  AO222X1 U109 ( .IN1(N489), .IN2(n93), .IN3(N209), .IN4(n94), .IN5(N197), 
        .IN6(n95), .Q(n125) );
  AO22X1 U110 ( .IN1(address[6]), .IN2(n493), .IN3(n84), .IN4(n126), .Q(n237)
         );
  OR2X1 U111 ( .IN1(n127), .IN2(n128), .Q(n126) );
  AO221X1 U112 ( .IN1(N146), .IN2(n503), .IN3(N113), .IN4(n501), .IN5(n129), 
        .Q(n128) );
  AO222X1 U113 ( .IN1(N370), .IN2(n509), .IN3(N124), .IN4(n89), .IN5(N359), 
        .IN6(n507), .Q(n129) );
  AO221X1 U114 ( .IN1(N478), .IN2(n90), .IN3(N314), .IN4(n91), .IN5(n130), .Q(
        n127) );
  AO222X1 U115 ( .IN1(N490), .IN2(n93), .IN3(N210), .IN4(n94), .IN5(N198), 
        .IN6(n95), .Q(n130) );
  AO22X1 U116 ( .IN1(n131), .IN2(n97), .IN3(address[7]), .IN4(n493), .Q(n238)
         );
  OR4X1 U117 ( .IN1(n132), .IN2(n133), .IN3(n134), .IN4(n135), .Q(n131) );
  AO222X1 U118 ( .IN1(N315), .IN2(n91), .IN3(N479), .IN4(n90), .IN5(N125), 
        .IN6(n89), .Q(n135) );
  AO222X1 U119 ( .IN1(N491), .IN2(n93), .IN3(N211), .IN4(n94), .IN5(N199), 
        .IN6(n95), .Q(n134) );
  AO21X1 U120 ( .IN1(N114), .IN2(n501), .IN3(n115), .Q(n133) );
  AO222X1 U121 ( .IN1(N360), .IN2(n507), .IN3(N371), .IN4(n509), .IN5(N147), 
        .IN6(n503), .Q(n132) );
  AO22X1 U122 ( .IN1(address[8]), .IN2(n493), .IN3(n84), .IN4(n136), .Q(n239)
         );
  OR2X1 U123 ( .IN1(n137), .IN2(n138), .Q(n136) );
  AO221X1 U124 ( .IN1(N148), .IN2(n503), .IN3(N115), .IN4(n501), .IN5(n139), 
        .Q(n138) );
  AO222X1 U125 ( .IN1(N372), .IN2(n509), .IN3(N126), .IN4(n89), .IN5(N361), 
        .IN6(n507), .Q(n139) );
  AO221X1 U126 ( .IN1(N480), .IN2(n90), .IN3(N316), .IN4(n91), .IN5(n140), .Q(
        n137) );
  AO222X1 U127 ( .IN1(N492), .IN2(n93), .IN3(N212), .IN4(n94), .IN5(N200), 
        .IN6(n95), .Q(n140) );
  AO22X1 U128 ( .IN1(n141), .IN2(n97), .IN3(address[9]), .IN4(n493), .Q(n240)
         );
  OR4X1 U129 ( .IN1(n142), .IN2(n143), .IN3(n144), .IN4(n145), .Q(n141) );
  AO222X1 U130 ( .IN1(N317), .IN2(n91), .IN3(N481), .IN4(n90), .IN5(N127), 
        .IN6(n89), .Q(n145) );
  AO222X1 U131 ( .IN1(N493), .IN2(n93), .IN3(N213), .IN4(n94), .IN5(N201), 
        .IN6(n95), .Q(n144) );
  AO21X1 U132 ( .IN1(N116), .IN2(n501), .IN3(n115), .Q(n143) );
  AO222X1 U133 ( .IN1(N362), .IN2(n507), .IN3(N373), .IN4(n509), .IN5(N149), 
        .IN6(n503), .Q(n142) );
  AO22X1 U134 ( .IN1(n146), .IN2(n97), .IN3(address[10]), .IN4(n493), .Q(n241)
         );
  NAND4X0 U135 ( .IN1(n147), .IN2(n148), .IN3(n499), .IN4(n149), .QN(n97) );
  NOR3X0 U136 ( .IN1(n150), .IN2(n509), .IN3(n151), .QN(n149) );
  OR4X1 U137 ( .IN1(n152), .IN2(n153), .IN3(n154), .IN4(n155), .Q(n146) );
  AO222X1 U138 ( .IN1(N318), .IN2(n91), .IN3(N482), .IN4(n90), .IN5(N128), 
        .IN6(n89), .Q(n155) );
  AO222X1 U139 ( .IN1(N494), .IN2(n93), .IN3(N214), .IN4(n94), .IN5(N202), 
        .IN6(n95), .Q(n154) );
  AO21X1 U140 ( .IN1(N117), .IN2(n501), .IN3(n115), .Q(n153) );
  AO222X1 U141 ( .IN1(N363), .IN2(n507), .IN3(N374), .IN4(n509), .IN5(N150), 
        .IN6(n503), .Q(n152) );
  AO22X1 U142 ( .IN1(k[15]), .IN2(n161), .IN3(N261), .IN4(n162), .Q(n242) );
  AO22X1 U143 ( .IN1(k[14]), .IN2(n161), .IN3(N260), .IN4(n162), .Q(n243) );
  AO22X1 U144 ( .IN1(k[13]), .IN2(n161), .IN3(N259), .IN4(n162), .Q(n244) );
  AO22X1 U145 ( .IN1(k[12]), .IN2(n161), .IN3(N258), .IN4(n162), .Q(n245) );
  AO22X1 U146 ( .IN1(k[11]), .IN2(n161), .IN3(N257), .IN4(n162), .Q(n246) );
  AO22X1 U147 ( .IN1(k[10]), .IN2(n161), .IN3(N256), .IN4(n162), .Q(n247) );
  AO22X1 U148 ( .IN1(k[9]), .IN2(n161), .IN3(N255), .IN4(n162), .Q(n248) );
  AO22X1 U149 ( .IN1(k[8]), .IN2(n161), .IN3(N254), .IN4(n162), .Q(n249) );
  AO22X1 U150 ( .IN1(k[7]), .IN2(n161), .IN3(N253), .IN4(n162), .Q(n250) );
  AO22X1 U151 ( .IN1(k[6]), .IN2(n161), .IN3(N252), .IN4(n162), .Q(n251) );
  AO22X1 U152 ( .IN1(k[5]), .IN2(n161), .IN3(N251), .IN4(n162), .Q(n252) );
  AO22X1 U153 ( .IN1(k[4]), .IN2(n161), .IN3(N250), .IN4(n162), .Q(n253) );
  AO22X1 U154 ( .IN1(k[3]), .IN2(n161), .IN3(N249), .IN4(n162), .Q(n254) );
  AO22X1 U155 ( .IN1(k[2]), .IN2(n161), .IN3(N248), .IN4(n162), .Q(n255) );
  AO22X1 U156 ( .IN1(N142), .IN2(n161), .IN3(N310), .IN4(n162), .Q(n256) );
  AO22X1 U157 ( .IN1(wr_en), .IN2(n494), .IN3(n163), .IN4(nrst), .Q(n257) );
  NAND4X0 U158 ( .IN1(n165), .IN2(n166), .IN3(n156), .IN4(n167), .QN(n164) );
  AO221X1 U159 ( .IN1(knownSinks[15]), .IN2(n168), .IN3(data_out[15]), .IN4(
        n169), .IN5(n170), .Q(n258) );
  AO22X1 U160 ( .IN1(N406), .IN2(n171), .IN3(N422), .IN4(n172), .Q(n170) );
  AO221X1 U161 ( .IN1(knownSinks[14]), .IN2(n168), .IN3(data_out[14]), .IN4(
        n169), .IN5(n173), .Q(n259) );
  AO22X1 U162 ( .IN1(N405), .IN2(n171), .IN3(N421), .IN4(n172), .Q(n173) );
  AO221X1 U163 ( .IN1(knownSinks[13]), .IN2(n168), .IN3(data_out[13]), .IN4(
        n169), .IN5(n174), .Q(n260) );
  AO22X1 U164 ( .IN1(N404), .IN2(n171), .IN3(N420), .IN4(n172), .Q(n174) );
  AO221X1 U165 ( .IN1(knownSinks[12]), .IN2(n168), .IN3(data_out[12]), .IN4(
        n169), .IN5(n175), .Q(n261) );
  AO22X1 U166 ( .IN1(N403), .IN2(n171), .IN3(N419), .IN4(n172), .Q(n175) );
  AO221X1 U167 ( .IN1(knownSinks[11]), .IN2(n168), .IN3(data_out[11]), .IN4(
        n169), .IN5(n176), .Q(n262) );
  AO22X1 U168 ( .IN1(N402), .IN2(n171), .IN3(N418), .IN4(n172), .Q(n176) );
  AO221X1 U169 ( .IN1(knownSinks[10]), .IN2(n168), .IN3(data_out[10]), .IN4(
        n169), .IN5(n177), .Q(n263) );
  AO22X1 U170 ( .IN1(N401), .IN2(n171), .IN3(N417), .IN4(n172), .Q(n177) );
  AO221X1 U171 ( .IN1(knownSinks[9]), .IN2(n168), .IN3(data_out[9]), .IN4(n169), .IN5(n178), .Q(n264) );
  AO22X1 U172 ( .IN1(N400), .IN2(n171), .IN3(N416), .IN4(n172), .Q(n178) );
  AO221X1 U173 ( .IN1(knownSinks[8]), .IN2(n168), .IN3(data_out[8]), .IN4(n169), .IN5(n179), .Q(n265) );
  AO22X1 U174 ( .IN1(N399), .IN2(n171), .IN3(N415), .IN4(n172), .Q(n179) );
  AO221X1 U175 ( .IN1(knownSinks[7]), .IN2(n168), .IN3(data_out[7]), .IN4(n169), .IN5(n180), .Q(n266) );
  AO22X1 U176 ( .IN1(N398), .IN2(n171), .IN3(N414), .IN4(n172), .Q(n180) );
  AO221X1 U177 ( .IN1(knownSinks[6]), .IN2(n168), .IN3(data_out[6]), .IN4(n169), .IN5(n181), .Q(n267) );
  AO22X1 U178 ( .IN1(N397), .IN2(n171), .IN3(N413), .IN4(n172), .Q(n181) );
  AO221X1 U179 ( .IN1(knownSinks[5]), .IN2(n168), .IN3(data_out[5]), .IN4(n169), .IN5(n182), .Q(n268) );
  AO22X1 U180 ( .IN1(N396), .IN2(n171), .IN3(N412), .IN4(n172), .Q(n182) );
  AO221X1 U181 ( .IN1(knownSinks[4]), .IN2(n168), .IN3(data_out[4]), .IN4(n169), .IN5(n183), .Q(n269) );
  AO22X1 U182 ( .IN1(N395), .IN2(n171), .IN3(N411), .IN4(n172), .Q(n183) );
  AO221X1 U183 ( .IN1(knownSinks[3]), .IN2(n168), .IN3(data_out[3]), .IN4(n169), .IN5(n184), .Q(n270) );
  AO22X1 U184 ( .IN1(N394), .IN2(n171), .IN3(N410), .IN4(n172), .Q(n184) );
  AO221X1 U185 ( .IN1(knownSinks[2]), .IN2(n168), .IN3(data_out[2]), .IN4(n169), .IN5(n185), .Q(n271) );
  AO22X1 U186 ( .IN1(N393), .IN2(n171), .IN3(N409), .IN4(n172), .Q(n185) );
  AO221X1 U187 ( .IN1(knownSinks[1]), .IN2(n168), .IN3(data_out[1]), .IN4(n169), .IN5(n186), .Q(n272) );
  AO22X1 U188 ( .IN1(N392), .IN2(n171), .IN3(N408), .IN4(n172), .Q(n186) );
  AO221X1 U189 ( .IN1(knownSinks[0]), .IN2(n168), .IN3(data_out[0]), .IN4(n169), .IN5(n187), .Q(n273) );
  AO22X1 U190 ( .IN1(N391), .IN2(n171), .IN3(N407), .IN4(n172), .Q(n187) );
  OR2X1 U191 ( .IN1(n492), .IN2(n169), .Q(n188) );
  AOI21X1 U193 ( .IN1(N262), .IN2(n91), .IN3(n505), .QN(n165) );
  AO22X1 U194 ( .IN1(j[14]), .IN2(n192), .IN3(N188), .IN4(n193), .Q(n274) );
  AO22X1 U195 ( .IN1(j[13]), .IN2(n192), .IN3(N187), .IN4(n193), .Q(n275) );
  AO22X1 U196 ( .IN1(j[12]), .IN2(n192), .IN3(N186), .IN4(n193), .Q(n276) );
  AO22X1 U197 ( .IN1(j[11]), .IN2(n192), .IN3(N185), .IN4(n193), .Q(n277) );
  AO22X1 U198 ( .IN1(j[10]), .IN2(n192), .IN3(N184), .IN4(n193), .Q(n278) );
  AO22X1 U199 ( .IN1(j[9]), .IN2(n192), .IN3(N183), .IN4(n193), .Q(n279) );
  AO22X1 U200 ( .IN1(j[8]), .IN2(n192), .IN3(N182), .IN4(n193), .Q(n280) );
  AO22X1 U201 ( .IN1(j[7]), .IN2(n192), .IN3(N181), .IN4(n193), .Q(n281) );
  AO22X1 U202 ( .IN1(j[6]), .IN2(n192), .IN3(N180), .IN4(n193), .Q(n282) );
  AO22X1 U203 ( .IN1(j[5]), .IN2(n192), .IN3(N179), .IN4(n193), .Q(n283) );
  AO22X1 U204 ( .IN1(j[4]), .IN2(n192), .IN3(N178), .IN4(n193), .Q(n284) );
  AO22X1 U205 ( .IN1(j[3]), .IN2(n192), .IN3(N177), .IN4(n193), .Q(n285) );
  AO22X1 U206 ( .IN1(j[2]), .IN2(n192), .IN3(N176), .IN4(n193), .Q(n286) );
  AO22X1 U207 ( .IN1(N109), .IN2(n192), .IN3(N194), .IN4(n193), .Q(n287) );
  AO22X1 U208 ( .IN1(N108), .IN2(n192), .IN3(N193), .IN4(n193), .Q(n288) );
  AO22X1 U209 ( .IN1(j[15]), .IN2(n192), .IN3(N189), .IN4(n193), .Q(n289) );
  AO22X1 U212 ( .IN1(i[15]), .IN2(n194), .IN3(N170), .IN4(n195), .Q(n290) );
  AO22X1 U213 ( .IN1(i[14]), .IN2(n194), .IN3(N169), .IN4(n195), .Q(n291) );
  AO22X1 U214 ( .IN1(i[13]), .IN2(n194), .IN3(N168), .IN4(n195), .Q(n292) );
  AO22X1 U215 ( .IN1(i[12]), .IN2(n194), .IN3(N167), .IN4(n195), .Q(n293) );
  AO22X1 U216 ( .IN1(i[11]), .IN2(n194), .IN3(N166), .IN4(n195), .Q(n294) );
  AO22X1 U217 ( .IN1(i[10]), .IN2(n194), .IN3(N165), .IN4(n195), .Q(n295) );
  AO22X1 U218 ( .IN1(i[9]), .IN2(n194), .IN3(N164), .IN4(n195), .Q(n296) );
  AO22X1 U219 ( .IN1(i[8]), .IN2(n194), .IN3(N163), .IN4(n195), .Q(n297) );
  AO22X1 U220 ( .IN1(i[7]), .IN2(n194), .IN3(N162), .IN4(n195), .Q(n298) );
  AO22X1 U221 ( .IN1(i[6]), .IN2(n194), .IN3(N161), .IN4(n195), .Q(n299) );
  AO22X1 U222 ( .IN1(i[5]), .IN2(n194), .IN3(N160), .IN4(n195), .Q(n300) );
  AO22X1 U223 ( .IN1(i[4]), .IN2(n194), .IN3(N159), .IN4(n195), .Q(n301) );
  AO22X1 U224 ( .IN1(i[3]), .IN2(n194), .IN3(N158), .IN4(n195), .Q(n302) );
  AO22X1 U225 ( .IN1(i[2]), .IN2(n194), .IN3(N157), .IN4(n195), .Q(n303) );
  AO22X1 U226 ( .IN1(N134), .IN2(n194), .IN3(N156), .IN4(n195), .Q(n304) );
  AO22X1 U227 ( .IN1(N133), .IN2(n194), .IN3(N155), .IN4(n195), .Q(n305) );
  AO22X1 U230 ( .IN1(neighborCount[15]), .IN2(n147), .IN3(data_in[15]), .IN4(
        n197), .Q(n306) );
  AO22X1 U231 ( .IN1(neighborCount[14]), .IN2(n147), .IN3(data_in[14]), .IN4(
        n197), .Q(n307) );
  AO22X1 U232 ( .IN1(neighborCount[13]), .IN2(n147), .IN3(data_in[13]), .IN4(
        n197), .Q(n308) );
  AO22X1 U233 ( .IN1(neighborCount[12]), .IN2(n147), .IN3(data_in[12]), .IN4(
        n197), .Q(n309) );
  AO22X1 U234 ( .IN1(neighborCount[11]), .IN2(n147), .IN3(data_in[11]), .IN4(
        n197), .Q(n310) );
  AO22X1 U235 ( .IN1(neighborCount[10]), .IN2(n147), .IN3(data_in[10]), .IN4(
        n197), .Q(n311) );
  AO22X1 U236 ( .IN1(neighborCount[9]), .IN2(n147), .IN3(data_in[9]), .IN4(
        n197), .Q(n312) );
  AO22X1 U237 ( .IN1(neighborCount[8]), .IN2(n147), .IN3(data_in[8]), .IN4(
        n197), .Q(n313) );
  AO22X1 U238 ( .IN1(neighborCount[7]), .IN2(n147), .IN3(data_in[7]), .IN4(
        n197), .Q(n314) );
  AO22X1 U239 ( .IN1(neighborCount[6]), .IN2(n147), .IN3(data_in[6]), .IN4(
        n197), .Q(n315) );
  AO22X1 U240 ( .IN1(neighborCount[5]), .IN2(n147), .IN3(data_in[5]), .IN4(
        n197), .Q(n316) );
  AO22X1 U241 ( .IN1(neighborCount[4]), .IN2(n147), .IN3(data_in[4]), .IN4(
        n197), .Q(n317) );
  AO22X1 U242 ( .IN1(neighborCount[3]), .IN2(n147), .IN3(data_in[3]), .IN4(
        n197), .Q(n318) );
  AO22X1 U243 ( .IN1(neighborCount[2]), .IN2(n147), .IN3(data_in[2]), .IN4(
        n197), .Q(n319) );
  AO22X1 U244 ( .IN1(neighborCount[1]), .IN2(n147), .IN3(data_in[1]), .IN4(
        n197), .Q(n320) );
  AO22X1 U245 ( .IN1(neighborCount[0]), .IN2(n147), .IN3(data_in[0]), .IN4(
        n197), .Q(n321) );
  AO22X1 U247 ( .IN1(knownSinkCount[15]), .IN2(n199), .IN3(n200), .IN4(
        data_in[15]), .Q(n322) );
  AO22X1 U248 ( .IN1(knownSinkCount[14]), .IN2(n199), .IN3(n200), .IN4(
        data_in[14]), .Q(n323) );
  AO22X1 U249 ( .IN1(knownSinkCount[13]), .IN2(n199), .IN3(n200), .IN4(
        data_in[13]), .Q(n324) );
  AO22X1 U250 ( .IN1(knownSinkCount[12]), .IN2(n199), .IN3(n200), .IN4(
        data_in[12]), .Q(n325) );
  AO22X1 U251 ( .IN1(knownSinkCount[11]), .IN2(n199), .IN3(n200), .IN4(
        data_in[11]), .Q(n326) );
  AO22X1 U252 ( .IN1(knownSinkCount[10]), .IN2(n199), .IN3(n200), .IN4(
        data_in[10]), .Q(n327) );
  AO22X1 U253 ( .IN1(knownSinkCount[9]), .IN2(n199), .IN3(n200), .IN4(
        data_in[9]), .Q(n328) );
  AO22X1 U254 ( .IN1(knownSinkCount[8]), .IN2(n199), .IN3(n200), .IN4(
        data_in[8]), .Q(n329) );
  AO22X1 U255 ( .IN1(knownSinkCount[7]), .IN2(n199), .IN3(n200), .IN4(
        data_in[7]), .Q(n330) );
  AO22X1 U256 ( .IN1(knownSinkCount[6]), .IN2(n199), .IN3(n200), .IN4(
        data_in[6]), .Q(n331) );
  AO22X1 U257 ( .IN1(knownSinkCount[5]), .IN2(n199), .IN3(n200), .IN4(
        data_in[5]), .Q(n332) );
  AO22X1 U258 ( .IN1(knownSinkCount[4]), .IN2(n199), .IN3(n200), .IN4(
        data_in[4]), .Q(n333) );
  AO22X1 U259 ( .IN1(knownSinkCount[3]), .IN2(n199), .IN3(n200), .IN4(
        data_in[3]), .Q(n334) );
  AO22X1 U260 ( .IN1(knownSinkCount[2]), .IN2(n199), .IN3(n200), .IN4(
        data_in[2]), .Q(n335) );
  AO22X1 U261 ( .IN1(knownSinkCount[1]), .IN2(n199), .IN3(n200), .IN4(
        data_in[1]), .Q(n336) );
  AO22X1 U262 ( .IN1(knownSinkCount[0]), .IN2(n199), .IN3(n200), .IN4(
        data_in[0]), .Q(n337) );
  AO22X1 U264 ( .IN1(n202), .IN2(knownSinks[15]), .IN3(n203), .IN4(data_in[15]), .Q(n338) );
  AO22X1 U265 ( .IN1(n202), .IN2(knownSinks[14]), .IN3(n203), .IN4(data_in[14]), .Q(n339) );
  AO22X1 U266 ( .IN1(n202), .IN2(knownSinks[13]), .IN3(n203), .IN4(data_in[13]), .Q(n340) );
  AO22X1 U267 ( .IN1(n202), .IN2(knownSinks[12]), .IN3(n203), .IN4(data_in[12]), .Q(n341) );
  AO22X1 U268 ( .IN1(n202), .IN2(knownSinks[11]), .IN3(n203), .IN4(data_in[11]), .Q(n342) );
  AO22X1 U269 ( .IN1(n202), .IN2(knownSinks[10]), .IN3(n203), .IN4(data_in[10]), .Q(n343) );
  AO22X1 U270 ( .IN1(n202), .IN2(knownSinks[9]), .IN3(n203), .IN4(data_in[9]), 
        .Q(n344) );
  AO22X1 U271 ( .IN1(n202), .IN2(knownSinks[8]), .IN3(n203), .IN4(data_in[8]), 
        .Q(n345) );
  AO22X1 U272 ( .IN1(n202), .IN2(knownSinks[7]), .IN3(n203), .IN4(data_in[7]), 
        .Q(n346) );
  AO22X1 U273 ( .IN1(n202), .IN2(knownSinks[6]), .IN3(n203), .IN4(data_in[6]), 
        .Q(n347) );
  AO22X1 U274 ( .IN1(n202), .IN2(knownSinks[5]), .IN3(n203), .IN4(data_in[5]), 
        .Q(n348) );
  AO22X1 U275 ( .IN1(n202), .IN2(knownSinks[4]), .IN3(n203), .IN4(data_in[4]), 
        .Q(n349) );
  AO22X1 U276 ( .IN1(n202), .IN2(knownSinks[3]), .IN3(n203), .IN4(data_in[3]), 
        .Q(n350) );
  AO22X1 U277 ( .IN1(n202), .IN2(knownSinks[2]), .IN3(n203), .IN4(data_in[2]), 
        .Q(n351) );
  AO22X1 U278 ( .IN1(n202), .IN2(knownSinks[1]), .IN3(n203), .IN4(data_in[1]), 
        .Q(n352) );
  AO22X1 U279 ( .IN1(n202), .IN2(knownSinks[0]), .IN3(n203), .IN4(data_in[0]), 
        .Q(n353) );
  AO22X1 U281 ( .IN1(done), .IN2(n166), .IN3(n508), .IN4(nrst), .Q(n354) );
  AO22X1 U282 ( .IN1(worstHops[15]), .IN2(n206), .IN3(n207), .IN4(data_in[15]), 
        .Q(n355) );
  AO22X1 U283 ( .IN1(worstHops[14]), .IN2(n206), .IN3(n207), .IN4(data_in[14]), 
        .Q(n356) );
  AO22X1 U284 ( .IN1(worstHops[13]), .IN2(n206), .IN3(n207), .IN4(data_in[13]), 
        .Q(n357) );
  AO22X1 U285 ( .IN1(worstHops[12]), .IN2(n206), .IN3(n207), .IN4(data_in[12]), 
        .Q(n358) );
  AO22X1 U286 ( .IN1(worstHops[11]), .IN2(n206), .IN3(n207), .IN4(data_in[11]), 
        .Q(n359) );
  AO22X1 U287 ( .IN1(worstHops[10]), .IN2(n206), .IN3(n207), .IN4(data_in[10]), 
        .Q(n360) );
  AO22X1 U288 ( .IN1(worstHops[9]), .IN2(n206), .IN3(n207), .IN4(data_in[9]), 
        .Q(n361) );
  AO22X1 U289 ( .IN1(worstHops[8]), .IN2(n206), .IN3(n207), .IN4(data_in[8]), 
        .Q(n362) );
  AO22X1 U290 ( .IN1(worstHops[7]), .IN2(n206), .IN3(n207), .IN4(data_in[7]), 
        .Q(n363) );
  AO22X1 U291 ( .IN1(worstHops[6]), .IN2(n206), .IN3(n207), .IN4(data_in[6]), 
        .Q(n364) );
  AO22X1 U292 ( .IN1(worstHops[5]), .IN2(n206), .IN3(n207), .IN4(data_in[5]), 
        .Q(n365) );
  AO22X1 U293 ( .IN1(worstHops[4]), .IN2(n206), .IN3(n207), .IN4(data_in[4]), 
        .Q(n366) );
  AO22X1 U294 ( .IN1(worstHops[3]), .IN2(n206), .IN3(n207), .IN4(data_in[3]), 
        .Q(n367) );
  AO22X1 U295 ( .IN1(worstHops[2]), .IN2(n206), .IN3(n207), .IN4(data_in[2]), 
        .Q(n368) );
  AO22X1 U296 ( .IN1(worstHops[1]), .IN2(n206), .IN3(n207), .IN4(data_in[1]), 
        .Q(n369) );
  AO22X1 U297 ( .IN1(worstHops[0]), .IN2(n206), .IN3(n207), .IN4(data_in[0]), 
        .Q(n370) );
  AO22X1 U299 ( .IN1(sinkIDCount[15]), .IN2(n208), .IN3(n209), .IN4(
        data_in[15]), .Q(n371) );
  AO22X1 U300 ( .IN1(sinkIDCount[14]), .IN2(n208), .IN3(n209), .IN4(
        data_in[14]), .Q(n372) );
  AO22X1 U301 ( .IN1(sinkIDCount[13]), .IN2(n208), .IN3(n209), .IN4(
        data_in[13]), .Q(n373) );
  AO22X1 U302 ( .IN1(sinkIDCount[12]), .IN2(n208), .IN3(n209), .IN4(
        data_in[12]), .Q(n374) );
  AO22X1 U303 ( .IN1(sinkIDCount[11]), .IN2(n208), .IN3(n209), .IN4(
        data_in[11]), .Q(n375) );
  AO22X1 U304 ( .IN1(sinkIDCount[10]), .IN2(n208), .IN3(n209), .IN4(
        data_in[10]), .Q(n376) );
  AO22X1 U305 ( .IN1(sinkIDCount[9]), .IN2(n208), .IN3(n209), .IN4(data_in[9]), 
        .Q(n377) );
  AO22X1 U306 ( .IN1(sinkIDCount[8]), .IN2(n208), .IN3(n209), .IN4(data_in[8]), 
        .Q(n378) );
  AO22X1 U307 ( .IN1(sinkIDCount[7]), .IN2(n208), .IN3(n209), .IN4(data_in[7]), 
        .Q(n379) );
  AO22X1 U308 ( .IN1(sinkIDCount[6]), .IN2(n208), .IN3(n209), .IN4(data_in[6]), 
        .Q(n380) );
  AO22X1 U309 ( .IN1(sinkIDCount[5]), .IN2(n208), .IN3(n209), .IN4(data_in[5]), 
        .Q(n381) );
  AO22X1 U310 ( .IN1(sinkIDCount[4]), .IN2(n208), .IN3(n209), .IN4(data_in[4]), 
        .Q(n382) );
  AO22X1 U311 ( .IN1(sinkIDCount[3]), .IN2(n208), .IN3(n209), .IN4(data_in[3]), 
        .Q(n383) );
  AO22X1 U312 ( .IN1(sinkIDCount[2]), .IN2(n208), .IN3(n209), .IN4(data_in[2]), 
        .Q(n384) );
  AO22X1 U313 ( .IN1(sinkIDCount[1]), .IN2(n208), .IN3(n209), .IN4(data_in[1]), 
        .Q(n385) );
  AO22X1 U314 ( .IN1(sinkIDCount[0]), .IN2(n208), .IN3(n209), .IN4(data_in[0]), 
        .Q(n386) );
  NAND4X0 U316 ( .IN1(n210), .IN2(n497), .IN3(n211), .IN4(n504), .QN(n387) );
  AO21X1 U317 ( .IN1(n212), .IN2(n510), .IN3(n91), .Q(n150) );
  NAND3X0 U319 ( .IN1(n198), .IN2(n189), .IN3(n216), .QN(n215) );
  NAND3X0 U320 ( .IN1(n190), .IN2(n498), .IN3(n148), .QN(n217) );
  AND3X1 U321 ( .IN1(n219), .IN2(n201), .IN3(n504), .Q(n148) );
  AND4X1 U322 ( .IN1(n196), .IN2(n158), .IN3(n222), .IN4(n223), .Q(n218) );
  NOR4X0 U323 ( .IN1(N262), .IN2(n501), .IN3(n220), .IN4(n89), .QN(n223) );
  NAND3X0 U324 ( .IN1(state[1]), .IN2(n71), .IN3(n224), .QN(n204) );
  NAND3X0 U325 ( .IN1(n225), .IN2(n81), .IN3(state[1]), .QN(n167) );
  AND3X1 U326 ( .IN1(n198), .IN2(n104), .IN3(n103), .Q(n158) );
  NAND3X0 U327 ( .IN1(n79), .IN2(n71), .IN3(n226), .QN(n104) );
  NAND3X0 U328 ( .IN1(n80), .IN2(n71), .IN3(n224), .QN(n198) );
  NAND4X0 U329 ( .IN1(n222), .IN2(n228), .IN3(n229), .IN4(n189), .QN(n389) );
  NAND3X0 U330 ( .IN1(n224), .IN2(n80), .IN3(state[3]), .QN(n189) );
  AND2X1 U331 ( .IN1(n156), .IN2(n157), .Q(n196) );
  OR2X1 U332 ( .IN1(n103), .IN2(en), .Q(n228) );
  AND3X1 U333 ( .IN1(n190), .IN2(n160), .IN3(n210), .Q(n222) );
  AND3X1 U334 ( .IN1(n230), .IN2(n205), .IN3(nrst), .Q(n210) );
  NAND3X0 U335 ( .IN1(n224), .IN2(state[1]), .IN3(state[3]), .QN(n205) );
  OR3X1 U336 ( .IN1(n79), .IN2(n226), .IN3(n71), .Q(n230) );
  NAND3X0 U337 ( .IN1(state[0]), .IN2(n225), .IN3(state[1]), .QN(n160) );
  NAND3X0 U338 ( .IN1(state[3]), .IN2(n79), .IN3(n226), .QN(n190) );
  AO22X1 U339 ( .IN1(N141), .IN2(n161), .IN3(N309), .IN4(n162), .Q(n390) );
  NAND3X0 U342 ( .IN1(state[3]), .IN2(state[2]), .IN3(n226), .QN(n103) );
  NOR3X0 U343 ( .IN1(state[0]), .IN2(state[2]), .IN3(n80), .QN(n227) );
  NAND3X0 U344 ( .IN1(n225), .IN2(n80), .IN3(state[0]), .QN(n191) );
  fixSinkList_DW01_inc_0 add_135 ( .A(sinkIDCount), .SUM({N422, N421, N420, 
        N419, N418, N417, N416, N415, N414, N413, N412, N411, N410, N409, N408, 
        N407}) );
  fixSinkList_DW01_inc_1 r235 ( .A({j[15:2], N109, N108}), .SUM({N189, N188, 
        N187, N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, 
        N194, N193}) );
  fixSinkList_DW01_inc_2 r233 ( .A({i[15:2], N134, N133}), .SUM({N170, N169, 
        N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, N158, N157, 
        N156, N155}) );
  fixSinkList_DW01_inc_3 add_96 ( .A({k[15:2], N142, N141}), .SUM({N261, N260, 
        N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, N248, 
        N310, N309}) );
  fixSinkList_DW01_inc_4 add_127 ( .A(worstHops), .SUM({N390, N389, N388, N387, 
        N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375}) );
  fixSinkList_DW01_add_11 add_127_2 ( .A(data_in), .B({N390, N389, N388, N387, 
        N386, N385, N384, N383, N382, N381, N380, N379, N378, N377, N376, N375}), .CI(1'b0), .SUM({N406, N405, N404, N403, N402, N401, N400, N399, N398, N397, 
        N396, N395, N394, N393, N392, N391}) );
  FADDX1 \add_0_root_add_67_2/U1_4  ( .A(k[3]), .B(N133), .CI(k[2]), .CO(
        \add_0_root_add_67_2/carry[5] ), .S(N144) );
  FADDX1 \add_0_root_add_67_2/U1_5  ( .A(k[4]), .B(N134), .CI(
        \add_0_root_add_67_2/carry[5] ), .CO(\add_0_root_add_67_2/carry[6] ), 
        .S(N145) );
  FADDX1 \add_0_root_add_67_2/U1_6  ( .A(k[5]), .B(N135), .CI(
        \add_0_root_add_67_2/carry[6] ), .CO(\add_0_root_add_67_2/carry[7] ), 
        .S(N146) );
  FADDX1 \add_0_root_add_67_2/U1_7  ( .A(k[6]), .B(N136), .CI(
        \add_0_root_add_67_2/carry[7] ), .CO(\add_0_root_add_67_2/carry[8] ), 
        .S(N147) );
  FADDX1 \add_0_root_add_67_2/U1_8  ( .A(k[7]), .B(N137), .CI(
        \add_0_root_add_67_2/carry[8] ), .CO(\add_0_root_add_67_2/carry[9] ), 
        .S(N148) );
  FADDX1 \add_0_root_add_67_2/U1_9  ( .A(k[8]), .B(N138), .CI(
        \add_0_root_add_67_2/carry[9] ), .CO(\add_0_root_add_67_2/carry[10] ), 
        .S(N149) );
  FADDX1 \add_0_root_add_67_2/U1_10  ( .A(k[9]), .B(N139), .CI(
        \add_0_root_add_67_2/carry[10] ), .S(N150) );
  FADDX1 \r241/U1_4  ( .A(N249), .B(N133), .CI(N248), .CO(\r241/carry[5] ), 
        .S(N312) );
  FADDX1 \r241/U1_5  ( .A(N250), .B(N134), .CI(\r241/carry[5] ), .CO(
        \r241/carry[6] ), .S(N313) );
  FADDX1 \r241/U1_6  ( .A(N251), .B(N135), .CI(\r241/carry[6] ), .CO(
        \r241/carry[7] ), .S(N314) );
  FADDX1 \r241/U1_7  ( .A(N252), .B(N136), .CI(\r241/carry[7] ), .CO(
        \r241/carry[8] ), .S(N315) );
  FADDX1 \r241/U1_8  ( .A(N253), .B(N137), .CI(\r241/carry[8] ), .CO(
        \r241/carry[9] ), .S(N316) );
  FADDX1 \r241/U1_9  ( .A(N254), .B(N138), .CI(\r241/carry[9] ), .CO(
        \r241/carry[10] ), .S(N317) );
  FADDX1 \r241/U1_10  ( .A(N255), .B(N139), .CI(\r241/carry[10] ), .S(N318) );
  DFFX1 done_buf_reg ( .D(n354), .CLK(clock), .Q(done) );
  DFFX1 \neighborCount_reg[15]  ( .D(n306), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n307), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n308), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n309), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n310), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n311), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n312), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n313), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n314), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n315), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n316), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n317), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n318), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n319), .CLK(clock), .Q(neighborCount[2])
         );
  DFFX1 \neighborCount_reg[1]  ( .D(n320), .CLK(clock), .Q(neighborCount[1]), 
        .QN(n466) );
  DFFX1 \neighborCount_reg[0]  ( .D(n321), .CLK(clock), .Q(neighborCount[0]), 
        .QN(n465) );
  DFFX1 \worstHops_reg[15]  ( .D(n355), .CLK(clock), .Q(worstHops[15]) );
  DFFX1 \worstHops_reg[14]  ( .D(n356), .CLK(clock), .Q(worstHops[14]) );
  DFFX1 \worstHops_reg[13]  ( .D(n357), .CLK(clock), .Q(worstHops[13]) );
  DFFX1 \worstHops_reg[12]  ( .D(n358), .CLK(clock), .Q(worstHops[12]) );
  DFFX1 \worstHops_reg[11]  ( .D(n359), .CLK(clock), .Q(worstHops[11]) );
  DFFX1 \worstHops_reg[10]  ( .D(n360), .CLK(clock), .Q(worstHops[10]) );
  DFFX1 \worstHops_reg[9]  ( .D(n361), .CLK(clock), .Q(worstHops[9]) );
  DFFX1 \worstHops_reg[8]  ( .D(n362), .CLK(clock), .Q(worstHops[8]) );
  DFFX1 \worstHops_reg[7]  ( .D(n363), .CLK(clock), .Q(worstHops[7]) );
  DFFX1 \worstHops_reg[6]  ( .D(n364), .CLK(clock), .Q(worstHops[6]) );
  DFFX1 \worstHops_reg[5]  ( .D(n365), .CLK(clock), .Q(worstHops[5]) );
  DFFX1 \worstHops_reg[4]  ( .D(n366), .CLK(clock), .Q(worstHops[4]) );
  DFFX1 \worstHops_reg[3]  ( .D(n367), .CLK(clock), .Q(worstHops[3]) );
  DFFX1 \worstHops_reg[2]  ( .D(n368), .CLK(clock), .Q(worstHops[2]) );
  DFFX1 \worstHops_reg[1]  ( .D(n369), .CLK(clock), .Q(worstHops[1]) );
  DFFX1 \worstHops_reg[0]  ( .D(n370), .CLK(clock), .Q(worstHops[0]) );
  DFFX1 \sinkIDCount_reg[15]  ( .D(n371), .CLK(clock), .Q(sinkIDCount[15]) );
  DFFX1 \sinkIDCount_reg[14]  ( .D(n372), .CLK(clock), .Q(sinkIDCount[14]) );
  DFFX1 \sinkIDCount_reg[13]  ( .D(n373), .CLK(clock), .Q(sinkIDCount[13]) );
  DFFX1 \sinkIDCount_reg[12]  ( .D(n374), .CLK(clock), .Q(sinkIDCount[12]) );
  DFFX1 \sinkIDCount_reg[11]  ( .D(n375), .CLK(clock), .Q(sinkIDCount[11]) );
  DFFX1 \sinkIDCount_reg[10]  ( .D(n376), .CLK(clock), .Q(sinkIDCount[10]) );
  DFFX1 \sinkIDCount_reg[9]  ( .D(n377), .CLK(clock), .Q(sinkIDCount[9]) );
  DFFX1 \sinkIDCount_reg[8]  ( .D(n378), .CLK(clock), .Q(sinkIDCount[8]) );
  DFFX1 \sinkIDCount_reg[7]  ( .D(n379), .CLK(clock), .Q(sinkIDCount[7]) );
  DFFX1 \sinkIDCount_reg[6]  ( .D(n380), .CLK(clock), .Q(sinkIDCount[6]) );
  DFFX1 \sinkIDCount_reg[5]  ( .D(n381), .CLK(clock), .Q(sinkIDCount[5]) );
  DFFX1 \sinkIDCount_reg[4]  ( .D(n382), .CLK(clock), .Q(sinkIDCount[4]) );
  DFFX1 \sinkIDCount_reg[3]  ( .D(n383), .CLK(clock), .Q(sinkIDCount[3]) );
  DFFX1 \sinkIDCount_reg[2]  ( .D(n384), .CLK(clock), .Q(sinkIDCount[2]) );
  DFFX1 \sinkIDCount_reg[1]  ( .D(n385), .CLK(clock), .Q(sinkIDCount[1]), .QN(
        n440) );
  DFFX1 \sinkIDCount_reg[0]  ( .D(n386), .CLK(clock), .Q(sinkIDCount[0]), .QN(
        n439) );
  DFFX1 \knownSinks_reg[15]  ( .D(n338), .CLK(clock), .Q(knownSinks[15]) );
  DFFX1 \knownSinks_reg[14]  ( .D(n339), .CLK(clock), .Q(knownSinks[14]) );
  DFFX1 \knownSinks_reg[13]  ( .D(n340), .CLK(clock), .Q(knownSinks[13]) );
  DFFX1 \knownSinks_reg[12]  ( .D(n341), .CLK(clock), .Q(knownSinks[12]) );
  DFFX1 \knownSinks_reg[11]  ( .D(n342), .CLK(clock), .Q(knownSinks[11]) );
  DFFX1 \knownSinks_reg[10]  ( .D(n343), .CLK(clock), .Q(knownSinks[10]) );
  DFFX1 \knownSinks_reg[9]  ( .D(n344), .CLK(clock), .Q(knownSinks[9]) );
  DFFX1 \knownSinks_reg[8]  ( .D(n345), .CLK(clock), .Q(knownSinks[8]) );
  DFFX1 \knownSinks_reg[7]  ( .D(n346), .CLK(clock), .Q(knownSinks[7]) );
  DFFX1 \knownSinks_reg[6]  ( .D(n347), .CLK(clock), .Q(knownSinks[6]) );
  DFFX1 \knownSinks_reg[5]  ( .D(n348), .CLK(clock), .Q(knownSinks[5]) );
  DFFX1 \knownSinks_reg[4]  ( .D(n349), .CLK(clock), .Q(knownSinks[4]) );
  DFFX1 \knownSinks_reg[3]  ( .D(n350), .CLK(clock), .Q(knownSinks[3]) );
  DFFX1 \knownSinks_reg[2]  ( .D(n351), .CLK(clock), .Q(knownSinks[2]) );
  DFFX1 \knownSinks_reg[1]  ( .D(n352), .CLK(clock), .Q(knownSinks[1]), .QN(
        n414) );
  DFFX1 \knownSinks_reg[0]  ( .D(n353), .CLK(clock), .Q(knownSinks[0]) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n322), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n323), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n324), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n325), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n326), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n327), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n328), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n329), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n330), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n331), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n332), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n333), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n334), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n335), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n336), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n491) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n337), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n490) );
  DFFX1 \k_reg[15]  ( .D(n242), .CLK(clock), .Q(k[15]) );
  DFFX1 \k_reg[14]  ( .D(n243), .CLK(clock), .Q(k[14]) );
  DFFX1 \k_reg[13]  ( .D(n244), .CLK(clock), .Q(k[13]) );
  DFFX1 \k_reg[12]  ( .D(n245), .CLK(clock), .Q(k[12]) );
  DFFX1 \k_reg[11]  ( .D(n246), .CLK(clock), .Q(k[11]) );
  DFFX1 \k_reg[10]  ( .D(n247), .CLK(clock), .Q(k[10]) );
  DFFX1 \k_reg[9]  ( .D(n248), .CLK(clock), .Q(k[9]) );
  DFFX1 \k_reg[8]  ( .D(n249), .CLK(clock), .Q(k[8]) );
  DFFX1 \k_reg[7]  ( .D(n250), .CLK(clock), .Q(k[7]) );
  DFFX1 \k_reg[6]  ( .D(n251), .CLK(clock), .Q(k[6]) );
  DFFX1 \k_reg[5]  ( .D(n252), .CLK(clock), .Q(k[5]) );
  DFFX1 \k_reg[4]  ( .D(n253), .CLK(clock), .Q(k[4]) );
  DFFX1 \k_reg[3]  ( .D(n254), .CLK(clock), .Q(k[3]) );
  DFFX1 \k_reg[2]  ( .D(n255), .CLK(clock), .Q(k[2]), .QN(N143) );
  DFFX1 \k_reg[1]  ( .D(n256), .CLK(clock), .Q(N142) );
  DFFX1 \k_reg[0]  ( .D(n390), .CLK(clock), .Q(N141) );
  DFFX1 wr_en_buf_reg ( .D(n257), .CLK(clock), .Q(wr_en) );
  DFFX1 \address_count_reg[0]  ( .D(n231), .CLK(clock), .Q(address[0]) );
  DFFX1 \i_reg[15]  ( .D(n290), .CLK(clock), .Q(i[15]) );
  DFFX1 \i_reg[14]  ( .D(n291), .CLK(clock), .Q(i[14]) );
  DFFX1 \i_reg[13]  ( .D(n292), .CLK(clock), .Q(i[13]) );
  DFFX1 \i_reg[12]  ( .D(n293), .CLK(clock), .Q(i[12]) );
  DFFX1 \i_reg[11]  ( .D(n294), .CLK(clock), .Q(i[11]) );
  DFFX1 \i_reg[10]  ( .D(n295), .CLK(clock), .Q(i[10]) );
  DFFX1 \i_reg[9]  ( .D(n296), .CLK(clock), .Q(i[9]) );
  DFFX1 \i_reg[8]  ( .D(n297), .CLK(clock), .Q(i[8]) );
  DFFX1 \i_reg[7]  ( .D(n298), .CLK(clock), .Q(i[7]) );
  DFFX1 \i_reg[6]  ( .D(n299), .CLK(clock), .Q(i[6]) );
  DFFX1 \i_reg[5]  ( .D(n300), .CLK(clock), .Q(i[5]) );
  DFFX1 \i_reg[4]  ( .D(n301), .CLK(clock), .Q(i[4]) );
  DFFX1 \i_reg[3]  ( .D(n302), .CLK(clock), .Q(i[3]) );
  DFFX1 \i_reg[2]  ( .D(n303), .CLK(clock), .Q(i[2]), .QN(N135) );
  DFFX1 \i_reg[1]  ( .D(n304), .CLK(clock), .Q(N134) );
  DFFX1 \i_reg[0]  ( .D(n305), .CLK(clock), .Q(N133), .QN(N119) );
  DFFX1 \address_count_reg[10]  ( .D(n241), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n240), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[7]  ( .D(n238), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[3]  ( .D(n234), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[1]  ( .D(n232), .CLK(clock), .Q(address[1]) );
  DFFX1 \j_reg[15]  ( .D(n289), .CLK(clock), .Q(j[15]) );
  DFFX1 \j_reg[14]  ( .D(n274), .CLK(clock), .Q(j[14]) );
  DFFX1 \j_reg[13]  ( .D(n275), .CLK(clock), .Q(j[13]) );
  DFFX1 \j_reg[12]  ( .D(n276), .CLK(clock), .Q(j[12]) );
  DFFX1 \j_reg[11]  ( .D(n277), .CLK(clock), .Q(j[11]) );
  DFFX1 \j_reg[10]  ( .D(n278), .CLK(clock), .Q(j[10]) );
  DFFX1 \j_reg[9]  ( .D(n279), .CLK(clock), .Q(j[9]) );
  DFFX1 \j_reg[8]  ( .D(n280), .CLK(clock), .Q(j[8]) );
  DFFX1 \j_reg[7]  ( .D(n281), .CLK(clock), .Q(j[7]) );
  DFFX1 \j_reg[6]  ( .D(n282), .CLK(clock), .Q(j[6]) );
  DFFX1 \j_reg[5]  ( .D(n283), .CLK(clock), .Q(j[5]) );
  DFFX1 \j_reg[4]  ( .D(n284), .CLK(clock), .Q(j[4]) );
  DFFX1 \j_reg[3]  ( .D(n285), .CLK(clock), .Q(j[3]) );
  DFFX1 \j_reg[2]  ( .D(n286), .CLK(clock), .Q(j[2]), .QN(N110) );
  DFFX1 \j_reg[1]  ( .D(n287), .CLK(clock), .Q(N109) );
  DFFX1 \j_reg[0]  ( .D(n288), .CLK(clock), .Q(N108) );
  DFFX1 \address_count_reg[8]  ( .D(n239), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[6]  ( .D(n237), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[5]  ( .D(n236), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n235), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[2]  ( .D(n233), .CLK(clock), .Q(address[2]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n265), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n266), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n267), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n268), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n269), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n270), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n271), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n272), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n273), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n264), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n263), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n262), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n261), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n260), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n259), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n258), .CLK(clock), .Q(data_out[15]) );
  NOR2X0 U345 ( .IN1(n510), .IN2(n157), .QN(n95) );
  INVX0 U346 ( .INP(n221), .ZN(n498) );
  INVX0 U347 ( .INP(n218), .ZN(n495) );
  NOR2X0 U348 ( .IN1(n157), .IN2(N171), .QN(n94) );
  NAND2X1 U349 ( .IN1(N152), .IN2(n502), .QN(n157) );
  INVX0 U350 ( .INP(n97), .ZN(n493) );
  NOR2X0 U351 ( .IN1(n510), .IN2(n196), .QN(n221) );
  INVX0 U352 ( .INP(N171), .ZN(n510) );
  NAND2X1 U353 ( .IN1(N171), .IN2(n212), .QN(n216) );
  INVX0 U354 ( .INP(n212), .ZN(n500) );
  INVX0 U355 ( .INP(n159), .ZN(n503) );
  INVX0 U356 ( .INP(n220), .ZN(n504) );
  NOR2X0 U357 ( .IN1(n191), .IN2(N152), .QN(n91) );
  NOR2X0 U358 ( .IN1(n188), .IN2(n189), .QN(n172) );
  NOR2X0 U359 ( .IN1(n190), .IN2(n188), .QN(n171) );
  INVX0 U360 ( .INP(n89), .ZN(n499) );
  NOR2X0 U361 ( .IN1(N190), .IN2(n500), .QN(n151) );
  NOR4X0 U362 ( .IN1(n492), .IN2(n194), .IN3(n500), .IN4(N171), .QN(n195) );
  NOR2X0 U363 ( .IN1(n188), .IN2(n191), .QN(n168) );
  NOR2X0 U364 ( .IN1(n204), .IN2(n492), .QN(n203) );
  NOR2X0 U365 ( .IN1(n160), .IN2(n492), .QN(n207) );
  NOR2X0 U366 ( .IN1(n198), .IN2(n492), .QN(n197) );
  NOR2X0 U367 ( .IN1(n201), .IN2(n492), .QN(n200) );
  NOR2X0 U368 ( .IN1(n159), .IN2(n492), .QN(n209) );
  AND2X1 U369 ( .IN1(n166), .IN2(n198), .Q(n147) );
  AND2X1 U370 ( .IN1(n166), .IN2(n498), .Q(n192) );
  AND2X1 U371 ( .IN1(n166), .IN2(n204), .Q(n202) );
  AND2X1 U372 ( .IN1(n166), .IN2(n160), .Q(n206) );
  AND2X1 U373 ( .IN1(n196), .IN2(n166), .Q(n194) );
  AND2X1 U374 ( .IN1(n166), .IN2(n201), .Q(n199) );
  AND2X1 U375 ( .IN1(n166), .IN2(n159), .Q(n208) );
  AND2X1 U376 ( .IN1(n500), .IN2(n166), .Q(n161) );
  NOR3X0 U377 ( .IN1(n192), .IN2(n500), .IN3(n492), .QN(n193) );
  NOR2X0 U378 ( .IN1(n492), .IN2(n493), .QN(n84) );
  INVX0 U379 ( .INP(N176), .ZN(N195) );
  NAND2X1 U380 ( .IN1(n103), .IN2(n104), .QN(n102) );
  INVX0 U381 ( .INP(N155), .ZN(N205) );
  NOR2X0 U382 ( .IN1(n492), .IN2(n218), .QN(n214) );
  AND2X1 U383 ( .IN1(n391), .IN2(n214), .Q(n388) );
  OR4X1 U384 ( .IN1(n215), .IN2(n507), .IN3(n91), .IN4(n501), .Q(n391) );
  NOR2X0 U385 ( .IN1(n156), .IN2(N171), .QN(n93) );
  NOR2X0 U386 ( .IN1(n510), .IN2(n156), .QN(n90) );
  INVX0 U387 ( .INP(N156), .ZN(n464) );
  INVX0 U388 ( .INP(N310), .ZN(n441) );
  NAND2X1 U389 ( .IN1(n226), .IN2(n225), .QN(n159) );
  NAND2X1 U390 ( .IN1(n204), .IN2(n189), .QN(n89) );
  INVX0 U391 ( .INP(n160), .ZN(n509) );
  NAND2X1 U392 ( .IN1(n191), .IN2(n156), .QN(n212) );
  INVX0 U393 ( .INP(n191), .ZN(n502) );
  INVX0 U394 ( .INP(n167), .ZN(n507) );
  NAND2X1 U395 ( .IN1(n159), .IN2(n167), .QN(n220) );
  INVX0 U396 ( .INP(n190), .ZN(n505) );
  INVX0 U397 ( .INP(n201), .ZN(n501) );
  INVX0 U398 ( .INP(N194), .ZN(n489) );
  AND3X1 U399 ( .IN1(nrst), .IN2(n189), .IN3(n165), .Q(n169) );
  INVX0 U400 ( .INP(data_in[1]), .ZN(n416) );
  INVX0 U401 ( .INP(data_in[0]), .ZN(n415) );
  NAND2X1 U402 ( .IN1(N190), .IN2(n221), .QN(n229) );
  AND2X1 U403 ( .IN1(n91), .IN2(nrst), .Q(n162) );
  OA21X1 U404 ( .IN1(en), .IN2(n103), .IN3(n204), .Q(n211) );
  INVX0 U405 ( .INP(n150), .ZN(n497) );
  OA21X1 U406 ( .IN1(n496), .IN2(n103), .IN3(nrst), .Q(n166) );
  INVX0 U407 ( .INP(en), .ZN(n496) );
  INVX0 U408 ( .INP(N248), .ZN(N311) );
  NAND2X1 U409 ( .IN1(start), .IN2(n506), .QN(n219) );
  INVX0 U410 ( .INP(n104), .ZN(n506) );
  NAND2X1 U411 ( .IN1(n158), .IN2(nrst), .QN(n115) );
  INVX0 U412 ( .INP(n164), .ZN(n494) );
  OA21X1 U413 ( .IN1(n505), .IN2(n502), .IN3(n164), .Q(n163) );
  INVX0 U414 ( .INP(n205), .ZN(n508) );
  INVX0 U415 ( .INP(nrst), .ZN(n492) );
  NOR2X0 U416 ( .IN1(n79), .IN2(state[3]), .QN(n225) );
  NAND2X1 U417 ( .IN1(n227), .IN2(n71), .QN(n201) );
  NAND2X1 U418 ( .IN1(n227), .IN2(state[3]), .QN(n156) );
  NOR2X0 U419 ( .IN1(state[1]), .IN2(state[0]), .QN(n226) );
  NOR2X0 U420 ( .IN1(n81), .IN2(state[2]), .QN(n224) );
  XNOR2X1 U421 ( .IN1(i[9]), .IN2(\r229/carry[10] ), .Q(N128) );
  OR2X1 U422 ( .IN1(i[8]), .IN2(\r229/carry[9] ), .Q(\r229/carry[10] ) );
  XNOR2X1 U423 ( .IN1(\r229/carry[9] ), .IN2(i[8]), .Q(N127) );
  AND2X1 U424 ( .IN1(\r229/carry[8] ), .IN2(i[7]), .Q(\r229/carry[9] ) );
  XOR2X1 U425 ( .IN1(i[7]), .IN2(\r229/carry[8] ), .Q(N126) );
  OR2X1 U426 ( .IN1(i[6]), .IN2(\r229/carry[7] ), .Q(\r229/carry[8] ) );
  XNOR2X1 U427 ( .IN1(\r229/carry[7] ), .IN2(i[6]), .Q(N125) );
  AND2X1 U428 ( .IN1(\r229/carry[6] ), .IN2(i[5]), .Q(\r229/carry[7] ) );
  XOR2X1 U429 ( .IN1(i[5]), .IN2(\r229/carry[6] ), .Q(N124) );
  AND2X1 U430 ( .IN1(\r229/carry[5] ), .IN2(i[4]), .Q(\r229/carry[6] ) );
  XOR2X1 U431 ( .IN1(i[4]), .IN2(\r229/carry[5] ), .Q(N123) );
  AND2X1 U432 ( .IN1(\r229/carry[4] ), .IN2(i[3]), .Q(\r229/carry[5] ) );
  XOR2X1 U433 ( .IN1(i[3]), .IN2(\r229/carry[4] ), .Q(N122) );
  OR2X1 U434 ( .IN1(i[2]), .IN2(\r229/carry[3] ), .Q(\r229/carry[4] ) );
  XNOR2X1 U435 ( .IN1(\r229/carry[3] ), .IN2(i[2]), .Q(N121) );
  OR2X1 U436 ( .IN1(N134), .IN2(N133), .Q(\r229/carry[3] ) );
  XNOR2X1 U437 ( .IN1(N133), .IN2(N134), .Q(N120) );
  XOR2X1 U438 ( .IN1(N183), .IN2(\add_155/carry[10] ), .Q(N482) );
  AND2X1 U439 ( .IN1(\add_155/carry[9] ), .IN2(N182), .Q(\add_155/carry[10] )
         );
  XOR2X1 U440 ( .IN1(N182), .IN2(\add_155/carry[9] ), .Q(N481) );
  AND2X1 U441 ( .IN1(\add_155/carry[8] ), .IN2(N181), .Q(\add_155/carry[9] )
         );
  XOR2X1 U442 ( .IN1(N181), .IN2(\add_155/carry[8] ), .Q(N480) );
  AND2X1 U443 ( .IN1(\add_155/carry[7] ), .IN2(N180), .Q(\add_155/carry[8] )
         );
  XOR2X1 U444 ( .IN1(N180), .IN2(\add_155/carry[7] ), .Q(N479) );
  AND2X1 U445 ( .IN1(\add_155/carry[6] ), .IN2(N179), .Q(\add_155/carry[7] )
         );
  XOR2X1 U446 ( .IN1(N179), .IN2(\add_155/carry[6] ), .Q(N478) );
  AND2X1 U447 ( .IN1(\add_155/carry[5] ), .IN2(N178), .Q(\add_155/carry[6] )
         );
  XOR2X1 U448 ( .IN1(N178), .IN2(\add_155/carry[5] ), .Q(N477) );
  AND2X1 U449 ( .IN1(N176), .IN2(N177), .Q(\add_155/carry[5] ) );
  XOR2X1 U450 ( .IN1(N177), .IN2(N176), .Q(N476) );
  XOR2X1 U451 ( .IN1(N183), .IN2(\add_87/carry[10] ), .Q(N202) );
  AND2X1 U452 ( .IN1(\add_87/carry[9] ), .IN2(N182), .Q(\add_87/carry[10] ) );
  XOR2X1 U453 ( .IN1(N182), .IN2(\add_87/carry[9] ), .Q(N201) );
  AND2X1 U454 ( .IN1(\add_87/carry[8] ), .IN2(N181), .Q(\add_87/carry[9] ) );
  XOR2X1 U455 ( .IN1(N181), .IN2(\add_87/carry[8] ), .Q(N200) );
  AND2X1 U456 ( .IN1(\add_87/carry[7] ), .IN2(N180), .Q(\add_87/carry[8] ) );
  XOR2X1 U457 ( .IN1(N180), .IN2(\add_87/carry[7] ), .Q(N199) );
  AND2X1 U458 ( .IN1(\add_87/carry[6] ), .IN2(N179), .Q(\add_87/carry[7] ) );
  XOR2X1 U459 ( .IN1(N179), .IN2(\add_87/carry[6] ), .Q(N198) );
  AND2X1 U460 ( .IN1(\add_87/carry[5] ), .IN2(N178), .Q(\add_87/carry[6] ) );
  XOR2X1 U461 ( .IN1(N178), .IN2(\add_87/carry[5] ), .Q(N197) );
  AND2X1 U462 ( .IN1(N176), .IN2(N177), .Q(\add_87/carry[5] ) );
  XOR2X1 U463 ( .IN1(N177), .IN2(N176), .Q(N196) );
  XNOR2X1 U464 ( .IN1(N164), .IN2(\add_92/carry[10] ), .Q(N214) );
  OR2X1 U465 ( .IN1(N163), .IN2(\add_92/carry[9] ), .Q(\add_92/carry[10] ) );
  XNOR2X1 U466 ( .IN1(\add_92/carry[9] ), .IN2(N163), .Q(N213) );
  AND2X1 U467 ( .IN1(\add_92/carry[8] ), .IN2(N162), .Q(\add_92/carry[9] ) );
  XOR2X1 U468 ( .IN1(N162), .IN2(\add_92/carry[8] ), .Q(N212) );
  OR2X1 U469 ( .IN1(N161), .IN2(\add_92/carry[7] ), .Q(\add_92/carry[8] ) );
  XNOR2X1 U470 ( .IN1(\add_92/carry[7] ), .IN2(N161), .Q(N211) );
  AND2X1 U471 ( .IN1(\add_92/carry[6] ), .IN2(N160), .Q(\add_92/carry[7] ) );
  XOR2X1 U472 ( .IN1(N160), .IN2(\add_92/carry[6] ), .Q(N210) );
  AND2X1 U473 ( .IN1(\add_92/carry[5] ), .IN2(N159), .Q(\add_92/carry[6] ) );
  XOR2X1 U474 ( .IN1(N159), .IN2(\add_92/carry[5] ), .Q(N209) );
  AND2X1 U475 ( .IN1(\add_92/carry[4] ), .IN2(N158), .Q(\add_92/carry[5] ) );
  XOR2X1 U476 ( .IN1(N158), .IN2(\add_92/carry[4] ), .Q(N208) );
  OR2X1 U477 ( .IN1(N157), .IN2(\add_92/carry[3] ), .Q(\add_92/carry[4] ) );
  XNOR2X1 U478 ( .IN1(\add_92/carry[3] ), .IN2(N157), .Q(N207) );
  OR2X1 U479 ( .IN1(N156), .IN2(N155), .Q(\add_92/carry[3] ) );
  XNOR2X1 U480 ( .IN1(N155), .IN2(N156), .Q(N206) );
  XNOR2X1 U481 ( .IN1(N164), .IN2(\add_160/carry[10] ), .Q(N494) );
  OR2X1 U482 ( .IN1(N163), .IN2(\add_160/carry[9] ), .Q(\add_160/carry[10] )
         );
  XNOR2X1 U483 ( .IN1(\add_160/carry[9] ), .IN2(N163), .Q(N493) );
  AND2X1 U484 ( .IN1(\add_160/carry[8] ), .IN2(N162), .Q(\add_160/carry[9] )
         );
  XOR2X1 U485 ( .IN1(N162), .IN2(\add_160/carry[8] ), .Q(N492) );
  OR2X1 U486 ( .IN1(N161), .IN2(\add_160/carry[7] ), .Q(\add_160/carry[8] ) );
  XNOR2X1 U487 ( .IN1(\add_160/carry[7] ), .IN2(N161), .Q(N491) );
  AND2X1 U488 ( .IN1(\add_160/carry[6] ), .IN2(N160), .Q(\add_160/carry[7] )
         );
  XOR2X1 U489 ( .IN1(N160), .IN2(\add_160/carry[6] ), .Q(N490) );
  AND2X1 U490 ( .IN1(\add_160/carry[5] ), .IN2(N159), .Q(\add_160/carry[6] )
         );
  XOR2X1 U491 ( .IN1(N159), .IN2(\add_160/carry[5] ), .Q(N489) );
  AND2X1 U492 ( .IN1(\add_160/carry[4] ), .IN2(N158), .Q(\add_160/carry[5] )
         );
  XOR2X1 U493 ( .IN1(N158), .IN2(\add_160/carry[4] ), .Q(N488) );
  OR2X1 U494 ( .IN1(N157), .IN2(\add_160/carry[3] ), .Q(\add_160/carry[4] ) );
  XNOR2X1 U495 ( .IN1(\add_160/carry[3] ), .IN2(N157), .Q(N487) );
  OR2X1 U496 ( .IN1(N156), .IN2(N155), .Q(\add_160/carry[3] ) );
  XNOR2X1 U497 ( .IN1(N155), .IN2(N156), .Q(N486) );
  XOR2X1 U498 ( .IN1(j[9]), .IN2(\add_55/carry[10] ), .Q(N117) );
  AND2X1 U499 ( .IN1(\add_55/carry[9] ), .IN2(j[8]), .Q(\add_55/carry[10] ) );
  XOR2X1 U500 ( .IN1(j[8]), .IN2(\add_55/carry[9] ), .Q(N116) );
  AND2X1 U501 ( .IN1(\add_55/carry[8] ), .IN2(j[7]), .Q(\add_55/carry[9] ) );
  XOR2X1 U502 ( .IN1(j[7]), .IN2(\add_55/carry[8] ), .Q(N115) );
  AND2X1 U503 ( .IN1(\add_55/carry[7] ), .IN2(j[6]), .Q(\add_55/carry[8] ) );
  XOR2X1 U504 ( .IN1(j[6]), .IN2(\add_55/carry[7] ), .Q(N114) );
  AND2X1 U505 ( .IN1(\add_55/carry[6] ), .IN2(j[5]), .Q(\add_55/carry[7] ) );
  XOR2X1 U506 ( .IN1(j[5]), .IN2(\add_55/carry[6] ), .Q(N113) );
  AND2X1 U507 ( .IN1(\add_55/carry[5] ), .IN2(j[4]), .Q(\add_55/carry[6] ) );
  XOR2X1 U508 ( .IN1(j[4]), .IN2(\add_55/carry[5] ), .Q(N112) );
  AND2X1 U509 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_55/carry[5] ) );
  XOR2X1 U510 ( .IN1(j[3]), .IN2(j[2]), .Q(N111) );
  XOR2X1 U511 ( .IN1(i[6]), .IN2(\r230/carry[10] ), .Q(N139) );
  OR2X1 U512 ( .IN1(i[5]), .IN2(\r230/carry[9] ), .Q(\r230/carry[10] ) );
  XNOR2X1 U513 ( .IN1(\r230/carry[9] ), .IN2(i[5]), .Q(N138) );
  AND2X1 U514 ( .IN1(\r230/carry[8] ), .IN2(i[4]), .Q(\r230/carry[9] ) );
  XOR2X1 U515 ( .IN1(i[4]), .IN2(\r230/carry[8] ), .Q(N137) );
  AND2X1 U516 ( .IN1(i[2]), .IN2(i[3]), .Q(\r230/carry[8] ) );
  XOR2X1 U517 ( .IN1(i[3]), .IN2(i[2]), .Q(N136) );
  XOR2X1 U518 ( .IN1(i[9]), .IN2(\add_121/carry[10] ), .Q(N374) );
  AND2X1 U519 ( .IN1(\add_121/carry[9] ), .IN2(i[8]), .Q(\add_121/carry[10] )
         );
  XOR2X1 U520 ( .IN1(i[8]), .IN2(\add_121/carry[9] ), .Q(N373) );
  OR2X1 U521 ( .IN1(i[7]), .IN2(\add_121/carry[8] ), .Q(\add_121/carry[9] ) );
  XNOR2X1 U522 ( .IN1(\add_121/carry[8] ), .IN2(i[7]), .Q(N372) );
  OR2X1 U523 ( .IN1(i[6]), .IN2(\add_121/carry[7] ), .Q(\add_121/carry[8] ) );
  XNOR2X1 U524 ( .IN1(\add_121/carry[7] ), .IN2(i[6]), .Q(N371) );
  OR2X1 U525 ( .IN1(i[5]), .IN2(\add_121/carry[6] ), .Q(\add_121/carry[7] ) );
  XNOR2X1 U526 ( .IN1(\add_121/carry[6] ), .IN2(i[5]), .Q(N370) );
  AND2X1 U527 ( .IN1(\add_121/carry[5] ), .IN2(i[4]), .Q(\add_121/carry[6] )
         );
  XOR2X1 U528 ( .IN1(i[4]), .IN2(\add_121/carry[5] ), .Q(N369) );
  AND2X1 U529 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_121/carry[5] ) );
  XOR2X1 U530 ( .IN1(i[3]), .IN2(i[2]), .Q(N368) );
  XOR2X1 U531 ( .IN1(j[9]), .IN2(\add_115/carry[10] ), .Q(N363) );
  AND2X1 U532 ( .IN1(\add_115/carry[9] ), .IN2(j[8]), .Q(\add_115/carry[10] )
         );
  XOR2X1 U533 ( .IN1(j[8]), .IN2(\add_115/carry[9] ), .Q(N362) );
  AND2X1 U534 ( .IN1(\add_115/carry[8] ), .IN2(j[7]), .Q(\add_115/carry[9] )
         );
  XOR2X1 U535 ( .IN1(j[7]), .IN2(\add_115/carry[8] ), .Q(N361) );
  AND2X1 U536 ( .IN1(\add_115/carry[7] ), .IN2(j[6]), .Q(\add_115/carry[8] )
         );
  XOR2X1 U537 ( .IN1(j[6]), .IN2(\add_115/carry[7] ), .Q(N360) );
  AND2X1 U538 ( .IN1(\add_115/carry[6] ), .IN2(j[5]), .Q(\add_115/carry[7] )
         );
  XOR2X1 U539 ( .IN1(j[5]), .IN2(\add_115/carry[6] ), .Q(N359) );
  OR2X1 U540 ( .IN1(j[4]), .IN2(\add_115/carry[5] ), .Q(\add_115/carry[6] ) );
  XNOR2X1 U541 ( .IN1(\add_115/carry[5] ), .IN2(j[4]), .Q(N358) );
  AND2X1 U542 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_115/carry[5] ) );
  XOR2X1 U543 ( .IN1(j[3]), .IN2(j[2]), .Q(N357) );
  XOR2X1 U544 ( .IN1(data_in[15]), .IN2(knownSinks[15]), .Q(n397) );
  XOR2X1 U545 ( .IN1(data_in[2]), .IN2(knownSinks[2]), .Q(n396) );
  NOR2X0 U546 ( .IN1(n415), .IN2(knownSinks[0]), .QN(n392) );
  OA22X1 U547 ( .IN1(data_in[1]), .IN2(n392), .IN3(n392), .IN4(n414), .Q(n395)
         );
  AND2X1 U548 ( .IN1(knownSinks[0]), .IN2(n415), .Q(n393) );
  OA22X1 U549 ( .IN1(n393), .IN2(n416), .IN3(knownSinks[1]), .IN4(n393), .Q(
        n394) );
  OR4X1 U550 ( .IN1(n397), .IN2(n396), .IN3(n395), .IN4(n394), .Q(n413) );
  XNOR2X1 U551 ( .IN1(data_in[6]), .IN2(knownSinks[6]), .Q(n401) );
  XNOR2X1 U552 ( .IN1(data_in[5]), .IN2(knownSinks[5]), .Q(n400) );
  XNOR2X1 U553 ( .IN1(data_in[4]), .IN2(knownSinks[4]), .Q(n399) );
  XNOR2X1 U554 ( .IN1(data_in[3]), .IN2(knownSinks[3]), .Q(n398) );
  NAND4X0 U555 ( .IN1(n401), .IN2(n400), .IN3(n399), .IN4(n398), .QN(n412) );
  XNOR2X1 U556 ( .IN1(data_in[10]), .IN2(knownSinks[10]), .Q(n405) );
  XNOR2X1 U557 ( .IN1(data_in[9]), .IN2(knownSinks[9]), .Q(n404) );
  XNOR2X1 U558 ( .IN1(data_in[8]), .IN2(knownSinks[8]), .Q(n403) );
  XNOR2X1 U559 ( .IN1(data_in[7]), .IN2(knownSinks[7]), .Q(n402) );
  NAND4X0 U560 ( .IN1(n405), .IN2(n404), .IN3(n403), .IN4(n402), .QN(n411) );
  XNOR2X1 U561 ( .IN1(data_in[14]), .IN2(knownSinks[14]), .Q(n409) );
  XNOR2X1 U562 ( .IN1(data_in[13]), .IN2(knownSinks[13]), .Q(n408) );
  XNOR2X1 U563 ( .IN1(data_in[12]), .IN2(knownSinks[12]), .Q(n407) );
  XNOR2X1 U564 ( .IN1(data_in[11]), .IN2(knownSinks[11]), .Q(n406) );
  NAND4X0 U565 ( .IN1(n409), .IN2(n408), .IN3(n407), .IN4(n406), .QN(n410) );
  NOR4X0 U566 ( .IN1(n413), .IN2(n412), .IN3(n411), .IN4(n410), .QN(N152) );
  XOR2X1 U567 ( .IN1(sinkIDCount[15]), .IN2(N261), .Q(n422) );
  XOR2X1 U568 ( .IN1(sinkIDCount[2]), .IN2(N248), .Q(n421) );
  NOR2X0 U569 ( .IN1(n439), .IN2(N309), .QN(n417) );
  OA22X1 U570 ( .IN1(sinkIDCount[1]), .IN2(n417), .IN3(n417), .IN4(n441), .Q(
        n420) );
  AND2X1 U571 ( .IN1(N309), .IN2(n439), .Q(n418) );
  OA22X1 U572 ( .IN1(n418), .IN2(n440), .IN3(N310), .IN4(n418), .Q(n419) );
  OR4X1 U573 ( .IN1(n422), .IN2(n421), .IN3(n420), .IN4(n419), .Q(n438) );
  XNOR2X1 U574 ( .IN1(sinkIDCount[6]), .IN2(N252), .Q(n426) );
  XNOR2X1 U575 ( .IN1(sinkIDCount[5]), .IN2(N251), .Q(n425) );
  XNOR2X1 U576 ( .IN1(sinkIDCount[4]), .IN2(N250), .Q(n424) );
  XNOR2X1 U577 ( .IN1(sinkIDCount[3]), .IN2(N249), .Q(n423) );
  NAND4X0 U578 ( .IN1(n426), .IN2(n425), .IN3(n424), .IN4(n423), .QN(n437) );
  XNOR2X1 U579 ( .IN1(sinkIDCount[10]), .IN2(N256), .Q(n430) );
  XNOR2X1 U580 ( .IN1(sinkIDCount[9]), .IN2(N255), .Q(n429) );
  XNOR2X1 U581 ( .IN1(sinkIDCount[8]), .IN2(N254), .Q(n428) );
  XNOR2X1 U582 ( .IN1(sinkIDCount[7]), .IN2(N253), .Q(n427) );
  NAND4X0 U583 ( .IN1(n430), .IN2(n429), .IN3(n428), .IN4(n427), .QN(n436) );
  XNOR2X1 U584 ( .IN1(sinkIDCount[14]), .IN2(N260), .Q(n434) );
  XNOR2X1 U585 ( .IN1(sinkIDCount[13]), .IN2(N259), .Q(n433) );
  XNOR2X1 U586 ( .IN1(sinkIDCount[12]), .IN2(N258), .Q(n432) );
  XNOR2X1 U587 ( .IN1(sinkIDCount[11]), .IN2(N257), .Q(n431) );
  NAND4X0 U588 ( .IN1(n434), .IN2(n433), .IN3(n432), .IN4(n431), .QN(n435) );
  NOR4X0 U589 ( .IN1(n438), .IN2(n437), .IN3(n436), .IN4(n435), .QN(N262) );
  XOR2X1 U590 ( .IN1(neighborCount[15]), .IN2(N170), .Q(n447) );
  XOR2X1 U591 ( .IN1(neighborCount[2]), .IN2(N157), .Q(n446) );
  NOR2X0 U592 ( .IN1(n465), .IN2(N155), .QN(n442) );
  OA22X1 U593 ( .IN1(neighborCount[1]), .IN2(n442), .IN3(n442), .IN4(n464), 
        .Q(n445) );
  AND2X1 U594 ( .IN1(N155), .IN2(n465), .Q(n443) );
  OA22X1 U595 ( .IN1(n443), .IN2(n466), .IN3(N156), .IN4(n443), .Q(n444) );
  OR4X1 U596 ( .IN1(n447), .IN2(n446), .IN3(n445), .IN4(n444), .Q(n463) );
  XNOR2X1 U597 ( .IN1(neighborCount[6]), .IN2(N161), .Q(n451) );
  XNOR2X1 U598 ( .IN1(neighborCount[5]), .IN2(N160), .Q(n450) );
  XNOR2X1 U599 ( .IN1(neighborCount[4]), .IN2(N159), .Q(n449) );
  XNOR2X1 U600 ( .IN1(neighborCount[3]), .IN2(N158), .Q(n448) );
  NAND4X0 U601 ( .IN1(n451), .IN2(n450), .IN3(n449), .IN4(n448), .QN(n462) );
  XNOR2X1 U602 ( .IN1(neighborCount[10]), .IN2(N165), .Q(n455) );
  XNOR2X1 U603 ( .IN1(neighborCount[9]), .IN2(N164), .Q(n454) );
  XNOR2X1 U604 ( .IN1(neighborCount[8]), .IN2(N163), .Q(n453) );
  XNOR2X1 U605 ( .IN1(neighborCount[7]), .IN2(N162), .Q(n452) );
  NAND4X0 U606 ( .IN1(n455), .IN2(n454), .IN3(n453), .IN4(n452), .QN(n461) );
  XNOR2X1 U607 ( .IN1(neighborCount[14]), .IN2(N169), .Q(n459) );
  XNOR2X1 U608 ( .IN1(neighborCount[13]), .IN2(N168), .Q(n458) );
  XNOR2X1 U609 ( .IN1(neighborCount[12]), .IN2(N167), .Q(n457) );
  XNOR2X1 U610 ( .IN1(neighborCount[11]), .IN2(N166), .Q(n456) );
  NAND4X0 U611 ( .IN1(n459), .IN2(n458), .IN3(n457), .IN4(n456), .QN(n460) );
  NOR4X0 U612 ( .IN1(n463), .IN2(n462), .IN3(n461), .IN4(n460), .QN(N171) );
  XOR2X1 U613 ( .IN1(knownSinkCount[15]), .IN2(N189), .Q(n472) );
  XOR2X1 U614 ( .IN1(knownSinkCount[2]), .IN2(N176), .Q(n471) );
  NOR2X0 U615 ( .IN1(n490), .IN2(N193), .QN(n467) );
  OA22X1 U616 ( .IN1(knownSinkCount[1]), .IN2(n467), .IN3(n467), .IN4(n489), 
        .Q(n470) );
  AND2X1 U617 ( .IN1(N193), .IN2(n490), .Q(n468) );
  OA22X1 U618 ( .IN1(n468), .IN2(n491), .IN3(N194), .IN4(n468), .Q(n469) );
  OR4X1 U619 ( .IN1(n472), .IN2(n471), .IN3(n470), .IN4(n469), .Q(n488) );
  XNOR2X1 U620 ( .IN1(knownSinkCount[6]), .IN2(N180), .Q(n476) );
  XNOR2X1 U621 ( .IN1(knownSinkCount[5]), .IN2(N179), .Q(n475) );
  XNOR2X1 U622 ( .IN1(knownSinkCount[4]), .IN2(N178), .Q(n474) );
  XNOR2X1 U623 ( .IN1(knownSinkCount[3]), .IN2(N177), .Q(n473) );
  NAND4X0 U624 ( .IN1(n476), .IN2(n475), .IN3(n474), .IN4(n473), .QN(n487) );
  XNOR2X1 U625 ( .IN1(knownSinkCount[10]), .IN2(N184), .Q(n480) );
  XNOR2X1 U626 ( .IN1(knownSinkCount[9]), .IN2(N183), .Q(n479) );
  XNOR2X1 U627 ( .IN1(knownSinkCount[8]), .IN2(N182), .Q(n478) );
  XNOR2X1 U628 ( .IN1(knownSinkCount[7]), .IN2(N181), .Q(n477) );
  NAND4X0 U629 ( .IN1(n480), .IN2(n479), .IN3(n478), .IN4(n477), .QN(n486) );
  XNOR2X1 U630 ( .IN1(knownSinkCount[14]), .IN2(N188), .Q(n484) );
  XNOR2X1 U631 ( .IN1(knownSinkCount[13]), .IN2(N187), .Q(n483) );
  XNOR2X1 U632 ( .IN1(knownSinkCount[12]), .IN2(N186), .Q(n482) );
  XNOR2X1 U633 ( .IN1(knownSinkCount[11]), .IN2(N185), .Q(n481) );
  NAND4X0 U634 ( .IN1(n484), .IN2(n483), .IN3(n482), .IN4(n481), .QN(n485) );
  NOR4X0 U635 ( .IN1(n488), .IN2(n487), .IN3(n486), .IN4(n485), .QN(N190) );
  AND2X1 U636 ( .IN1(address[0]), .IN2(n493), .Q(n231) );
endmodule

