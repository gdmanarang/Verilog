
module neighborSinkInOtherCluster_DW01_inc_0 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module neighborSinkInOtherCluster_DW01_inc_1 ( A, SUM );
  input [15:0] A;
  output [15:0] SUM;

  wire   [15:2] carry;

  HADDX1 U1_1_14 ( .A0(A[14]), .B0(carry[14]), .C1(carry[15]), .SO(SUM[14]) );
  HADDX1 U1_1_13 ( .A0(A[13]), .B0(carry[13]), .C1(carry[14]), .SO(SUM[13]) );
  HADDX1 U1_1_12 ( .A0(A[12]), .B0(carry[12]), .C1(carry[13]), .SO(SUM[12]) );
  HADDX1 U1_1_11 ( .A0(A[11]), .B0(carry[11]), .C1(carry[12]), .SO(SUM[11]) );
  HADDX1 U1_1_10 ( .A0(A[10]), .B0(carry[10]), .C1(carry[11]), .SO(SUM[10]) );
  HADDX1 U1_1_9 ( .A0(A[9]), .B0(carry[9]), .C1(carry[10]), .SO(SUM[9]) );
  HADDX1 U1_1_8 ( .A0(A[8]), .B0(carry[8]), .C1(carry[9]), .SO(SUM[8]) );
  HADDX1 U1_1_7 ( .A0(A[7]), .B0(carry[7]), .C1(carry[8]), .SO(SUM[7]) );
  HADDX1 U1_1_6 ( .A0(A[6]), .B0(carry[6]), .C1(carry[7]), .SO(SUM[6]) );
  HADDX1 U1_1_5 ( .A0(A[5]), .B0(carry[5]), .C1(carry[6]), .SO(SUM[5]) );
  HADDX1 U1_1_4 ( .A0(A[4]), .B0(carry[4]), .C1(carry[5]), .SO(SUM[4]) );
  HADDX1 U1_1_3 ( .A0(A[3]), .B0(carry[3]), .C1(carry[4]), .SO(SUM[3]) );
  HADDX1 U1_1_2 ( .A0(A[2]), .B0(carry[2]), .C1(carry[3]), .SO(SUM[2]) );
  HADDX1 U1_1_1 ( .A0(A[1]), .B0(A[0]), .C1(carry[2]), .SO(SUM[1]) );
  INVX0 U1 ( .INP(A[0]), .ZN(SUM[0]) );
  XOR2X1 U2 ( .IN1(carry[15]), .IN2(A[15]), .Q(SUM[15]) );
endmodule


module neighborSinkInOtherCluster ( clock, nrst, en, start, address, wr_en, 
        data_in, MY_CLUSTER_ID, data_out, forAggregation, done );
  output [10:0] address;
  input [15:0] data_in;
  input [15:0] MY_CLUSTER_ID;
  output [15:0] data_out;
  input clock, nrst, en, start;
  output wr_en, forAggregation, done;
  wire   N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N91, N92, N93, N94,
         N95, N96, N97, N98, N99, N100, N102, N103, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N136,
         N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
         N148, N149, N151, N152, N153, N154, N155, N156, N157, N158, N159,
         N160, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, n23, n29, n30, n31, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, \add_92/carry[10] , \add_92/carry[9] ,
         \add_92/carry[8] , \add_92/carry[7] , \add_92/carry[6] ,
         \add_92/carry[5] , \add_86/carry[10] , \add_86/carry[9] ,
         \add_86/carry[8] , \add_86/carry[7] , \add_86/carry[6] ,
         \add_86/carry[5] , \add_72/carry[10] , \add_72/carry[9] ,
         \add_72/carry[8] , \add_72/carry[7] , \add_72/carry[6] ,
         \add_72/carry[5] , \add_66/carry[10] , \add_66/carry[9] ,
         \add_66/carry[8] , \add_66/carry[7] , \add_66/carry[6] ,
         \add_66/carry[5] , n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337;
  wire   [3:0] state;
  wire   [15:0] i;
  wire   [15:0] j;
  wire   [15:0] clusterID;
  wire   [15:0] knownSinkCount;
  wire   [15:0] neighborCount;
  wire   [15:0] neighborID;
  assign data_out[15] = 1'b0;
  assign data_out[14] = 1'b0;
  assign data_out[13] = 1'b0;
  assign data_out[12] = 1'b0;
  assign data_out[11] = 1'b0;
  assign data_out[10] = 1'b0;
  assign data_out[9] = 1'b0;
  assign data_out[8] = 1'b0;
  assign data_out[7] = 1'b0;
  assign data_out[6] = 1'b0;
  assign data_out[5] = 1'b0;
  assign data_out[4] = 1'b0;
  assign data_out[3] = 1'b0;
  assign data_out[2] = 1'b0;
  assign data_out[1] = 1'b0;

  DFFX1 \state_reg[0]  ( .D(n218), .CLK(clock), .Q(state[0]), .QN(n31) );
  DFFX1 \state_reg[2]  ( .D(n216), .CLK(clock), .Q(state[2]), .QN(n29) );
  DFFX1 \state_reg[1]  ( .D(n217), .CLK(clock), .Q(state[1]), .QN(n30) );
  DFFX1 \state_reg[3]  ( .D(n219), .CLK(clock), .Q(state[3]), .QN(n23) );
  AO22X1 U69 ( .IN1(wr_en), .IN2(n330), .IN3(n36), .IN4(n37), .Q(n106) );
  NAND3X0 U70 ( .IN1(n38), .IN2(n39), .IN3(n40), .QN(n37) );
  AO22X1 U71 ( .IN1(done), .IN2(n325), .IN3(n334), .IN4(nrst), .Q(n107) );
  AO22X1 U72 ( .IN1(forAggregation), .IN2(n42), .IN3(n36), .IN4(n332), .Q(n108) );
  AO22X1 U73 ( .IN1(n43), .IN2(n44), .IN3(address[10]), .IN4(n324), .Q(n109)
         );
  AO221X1 U74 ( .IN1(n45), .IN2(n46), .IN3(N100), .IN4(n337), .IN5(n47), .Q(
        n44) );
  AO21X1 U75 ( .IN1(N89), .IN2(n333), .IN3(n326), .Q(n47) );
  AO22X1 U76 ( .IN1(N160), .IN2(n222), .IN3(N131), .IN4(n223), .Q(n46) );
  AO22X1 U77 ( .IN1(n48), .IN2(n43), .IN3(address[9]), .IN4(n324), .Q(n110) );
  AO221X1 U78 ( .IN1(n45), .IN2(n49), .IN3(N99), .IN4(n337), .IN5(n50), .Q(n48) );
  AO21X1 U79 ( .IN1(N88), .IN2(n333), .IN3(n326), .Q(n50) );
  AO22X1 U80 ( .IN1(N159), .IN2(n222), .IN3(N130), .IN4(n223), .Q(n49) );
  AO221X1 U81 ( .IN1(N158), .IN2(n51), .IN3(address[8]), .IN4(n324), .IN5(n52), 
        .Q(n111) );
  AO222X1 U82 ( .IN1(N87), .IN2(n53), .IN3(N98), .IN4(n54), .IN5(N129), .IN6(
        n55), .Q(n52) );
  AO22X1 U83 ( .IN1(n56), .IN2(n43), .IN3(address[7]), .IN4(n324), .Q(n112) );
  AO221X1 U84 ( .IN1(n45), .IN2(n57), .IN3(N97), .IN4(n337), .IN5(n58), .Q(n56) );
  AO21X1 U85 ( .IN1(N86), .IN2(n333), .IN3(n326), .Q(n58) );
  AO22X1 U86 ( .IN1(N157), .IN2(n222), .IN3(N128), .IN4(n223), .Q(n57) );
  AO221X1 U87 ( .IN1(nrst), .IN2(n60), .IN3(address[6]), .IN4(n324), .IN5(n61), 
        .Q(n113) );
  AO22X1 U88 ( .IN1(N156), .IN2(n51), .IN3(N127), .IN4(n55), .Q(n61) );
  AO221X1 U89 ( .IN1(N96), .IN2(n337), .IN3(N85), .IN4(n333), .IN5(n336), .Q(
        n60) );
  AO221X1 U90 ( .IN1(N155), .IN2(n51), .IN3(address[5]), .IN4(n324), .IN5(n62), 
        .Q(n114) );
  AO222X1 U91 ( .IN1(N84), .IN2(n53), .IN3(N95), .IN4(n54), .IN5(N126), .IN6(
        n55), .Q(n62) );
  AO221X1 U92 ( .IN1(N154), .IN2(n51), .IN3(address[4]), .IN4(n324), .IN5(n63), 
        .Q(n115) );
  AO222X1 U93 ( .IN1(N83), .IN2(n53), .IN3(N94), .IN4(n54), .IN5(N125), .IN6(
        n55), .Q(n63) );
  AO22X1 U94 ( .IN1(n64), .IN2(n43), .IN3(address[3]), .IN4(n324), .Q(n116) );
  NAND3X0 U95 ( .IN1(n59), .IN2(n65), .IN3(n66), .QN(n64) );
  AOI221X1 U96 ( .IN1(N93), .IN2(n337), .IN3(n45), .IN4(n67), .IN5(n336), .QN(
        n66) );
  AO22X1 U97 ( .IN1(N153), .IN2(n222), .IN3(N124), .IN4(n223), .Q(n67) );
  NOR4X0 U98 ( .IN1(n328), .IN2(n335), .IN3(n41), .IN4(n69), .QN(n59) );
  AO221X1 U99 ( .IN1(N152), .IN2(n51), .IN3(address[2]), .IN4(n324), .IN5(n70), 
        .Q(n117) );
  AO222X1 U100 ( .IN1(N81), .IN2(n53), .IN3(N92), .IN4(n54), .IN5(N123), .IN6(
        n55), .Q(n70) );
  AO222X1 U101 ( .IN1(nrst), .IN2(n71), .IN3(n36), .IN4(n72), .IN5(address[1]), 
        .IN6(n324), .Q(n118) );
  AO221X1 U102 ( .IN1(N122), .IN2(n223), .IN3(N151), .IN4(n222), .IN5(n332), 
        .Q(n72) );
  AO221X1 U103 ( .IN1(N91), .IN2(n337), .IN3(N80), .IN4(n333), .IN5(n335), .Q(
        n71) );
  AND2X1 U106 ( .IN1(n74), .IN2(n223), .Q(n55) );
  NAND4X0 U107 ( .IN1(n75), .IN2(n42), .IN3(n76), .IN4(n77), .QN(n43) );
  AND2X1 U108 ( .IN1(n74), .IN2(n222), .Q(n51) );
  AO22X1 U109 ( .IN1(nrst), .IN2(n329), .IN3(data_out[0]), .IN4(n39), .Q(n120)
         );
  AO22X1 U110 ( .IN1(i[14]), .IN2(n78), .IN3(N148), .IN4(n79), .Q(n121) );
  AO22X1 U111 ( .IN1(i[13]), .IN2(n78), .IN3(N147), .IN4(n79), .Q(n122) );
  AO22X1 U112 ( .IN1(i[12]), .IN2(n78), .IN3(N146), .IN4(n79), .Q(n123) );
  AO22X1 U113 ( .IN1(i[11]), .IN2(n78), .IN3(N145), .IN4(n79), .Q(n124) );
  AO22X1 U114 ( .IN1(i[10]), .IN2(n78), .IN3(N144), .IN4(n79), .Q(n125) );
  AO22X1 U115 ( .IN1(i[9]), .IN2(n78), .IN3(N143), .IN4(n79), .Q(n126) );
  AO22X1 U116 ( .IN1(i[8]), .IN2(n78), .IN3(N142), .IN4(n79), .Q(n127) );
  AO22X1 U117 ( .IN1(i[7]), .IN2(n78), .IN3(N141), .IN4(n79), .Q(n128) );
  AO22X1 U118 ( .IN1(i[6]), .IN2(n78), .IN3(N140), .IN4(n79), .Q(n129) );
  AO22X1 U119 ( .IN1(i[5]), .IN2(n78), .IN3(N139), .IN4(n79), .Q(n130) );
  AO22X1 U120 ( .IN1(i[4]), .IN2(n78), .IN3(N138), .IN4(n79), .Q(n131) );
  AO22X1 U121 ( .IN1(i[3]), .IN2(n78), .IN3(N137), .IN4(n79), .Q(n132) );
  AO22X1 U122 ( .IN1(i[2]), .IN2(n78), .IN3(N136), .IN4(n79), .Q(n133) );
  AO22X1 U123 ( .IN1(N81), .IN2(n78), .IN3(N152), .IN4(n79), .Q(n134) );
  AO22X1 U124 ( .IN1(N80), .IN2(n78), .IN3(N151), .IN4(n79), .Q(n135) );
  AO22X1 U125 ( .IN1(i[15]), .IN2(n78), .IN3(N149), .IN4(n79), .Q(n136) );
  AO22X1 U126 ( .IN1(j[15]), .IN2(n42), .IN3(N120), .IN4(n80), .Q(n137) );
  AO22X1 U127 ( .IN1(j[14]), .IN2(n42), .IN3(N119), .IN4(n80), .Q(n138) );
  AO22X1 U128 ( .IN1(j[13]), .IN2(n42), .IN3(N118), .IN4(n80), .Q(n139) );
  AO22X1 U129 ( .IN1(j[12]), .IN2(n42), .IN3(N117), .IN4(n80), .Q(n140) );
  AO22X1 U130 ( .IN1(j[11]), .IN2(n42), .IN3(N116), .IN4(n80), .Q(n141) );
  AO22X1 U131 ( .IN1(j[10]), .IN2(n42), .IN3(N115), .IN4(n80), .Q(n142) );
  AO22X1 U132 ( .IN1(j[9]), .IN2(n42), .IN3(N114), .IN4(n80), .Q(n143) );
  AO22X1 U133 ( .IN1(j[8]), .IN2(n42), .IN3(N113), .IN4(n80), .Q(n144) );
  AO22X1 U134 ( .IN1(j[7]), .IN2(n42), .IN3(N112), .IN4(n80), .Q(n145) );
  AO22X1 U135 ( .IN1(j[6]), .IN2(n42), .IN3(N111), .IN4(n80), .Q(n146) );
  AO22X1 U136 ( .IN1(j[5]), .IN2(n42), .IN3(N110), .IN4(n80), .Q(n147) );
  AO22X1 U137 ( .IN1(j[4]), .IN2(n42), .IN3(N109), .IN4(n80), .Q(n148) );
  AO22X1 U138 ( .IN1(j[3]), .IN2(n42), .IN3(N108), .IN4(n80), .Q(n149) );
  AO22X1 U139 ( .IN1(j[2]), .IN2(n42), .IN3(N107), .IN4(n80), .Q(n150) );
  AO22X1 U140 ( .IN1(N92), .IN2(n42), .IN3(N123), .IN4(n80), .Q(n151) );
  AO22X1 U141 ( .IN1(N91), .IN2(n42), .IN3(N122), .IN4(n80), .Q(n152) );
  AO22X1 U143 ( .IN1(knownSinkCount[15]), .IN2(n82), .IN3(data_in[15]), .IN4(
        n83), .Q(n153) );
  AO22X1 U144 ( .IN1(knownSinkCount[14]), .IN2(n82), .IN3(data_in[14]), .IN4(
        n83), .Q(n154) );
  AO22X1 U145 ( .IN1(knownSinkCount[13]), .IN2(n82), .IN3(data_in[13]), .IN4(
        n83), .Q(n155) );
  AO22X1 U146 ( .IN1(knownSinkCount[12]), .IN2(n82), .IN3(data_in[12]), .IN4(
        n83), .Q(n156) );
  AO22X1 U147 ( .IN1(knownSinkCount[11]), .IN2(n82), .IN3(data_in[11]), .IN4(
        n83), .Q(n157) );
  AO22X1 U148 ( .IN1(knownSinkCount[10]), .IN2(n82), .IN3(data_in[10]), .IN4(
        n83), .Q(n158) );
  AO22X1 U149 ( .IN1(knownSinkCount[9]), .IN2(n82), .IN3(data_in[9]), .IN4(n83), .Q(n159) );
  AO22X1 U150 ( .IN1(knownSinkCount[8]), .IN2(n82), .IN3(data_in[8]), .IN4(n83), .Q(n160) );
  AO22X1 U151 ( .IN1(knownSinkCount[7]), .IN2(n82), .IN3(data_in[7]), .IN4(n83), .Q(n161) );
  AO22X1 U152 ( .IN1(knownSinkCount[6]), .IN2(n82), .IN3(data_in[6]), .IN4(n83), .Q(n162) );
  AO22X1 U153 ( .IN1(knownSinkCount[5]), .IN2(n82), .IN3(data_in[5]), .IN4(n83), .Q(n163) );
  AO22X1 U154 ( .IN1(knownSinkCount[4]), .IN2(n82), .IN3(data_in[4]), .IN4(n83), .Q(n164) );
  AO22X1 U155 ( .IN1(knownSinkCount[3]), .IN2(n82), .IN3(data_in[3]), .IN4(n83), .Q(n165) );
  AO22X1 U156 ( .IN1(knownSinkCount[2]), .IN2(n82), .IN3(data_in[2]), .IN4(n83), .Q(n166) );
  AO22X1 U157 ( .IN1(knownSinkCount[1]), .IN2(n82), .IN3(data_in[1]), .IN4(n83), .Q(n167) );
  AO22X1 U158 ( .IN1(knownSinkCount[0]), .IN2(n82), .IN3(data_in[0]), .IN4(n83), .Q(n168) );
  AO22X1 U159 ( .IN1(neighborCount[15]), .IN2(n84), .IN3(n85), .IN4(
        data_in[15]), .Q(n169) );
  AO22X1 U160 ( .IN1(neighborCount[14]), .IN2(n84), .IN3(n85), .IN4(
        data_in[14]), .Q(n170) );
  AO22X1 U161 ( .IN1(neighborCount[13]), .IN2(n84), .IN3(n85), .IN4(
        data_in[13]), .Q(n171) );
  AO22X1 U162 ( .IN1(neighborCount[12]), .IN2(n84), .IN3(n85), .IN4(
        data_in[12]), .Q(n172) );
  AO22X1 U163 ( .IN1(neighborCount[11]), .IN2(n84), .IN3(n85), .IN4(
        data_in[11]), .Q(n173) );
  AO22X1 U164 ( .IN1(neighborCount[10]), .IN2(n84), .IN3(n85), .IN4(
        data_in[10]), .Q(n174) );
  AO22X1 U165 ( .IN1(neighborCount[9]), .IN2(n84), .IN3(n85), .IN4(data_in[9]), 
        .Q(n175) );
  AO22X1 U166 ( .IN1(neighborCount[8]), .IN2(n84), .IN3(n85), .IN4(data_in[8]), 
        .Q(n176) );
  AO22X1 U167 ( .IN1(neighborCount[7]), .IN2(n84), .IN3(n85), .IN4(data_in[7]), 
        .Q(n177) );
  AO22X1 U168 ( .IN1(neighborCount[6]), .IN2(n84), .IN3(n85), .IN4(data_in[6]), 
        .Q(n178) );
  AO22X1 U169 ( .IN1(neighborCount[5]), .IN2(n84), .IN3(n85), .IN4(data_in[5]), 
        .Q(n179) );
  AO22X1 U170 ( .IN1(neighborCount[4]), .IN2(n84), .IN3(n85), .IN4(data_in[4]), 
        .Q(n180) );
  AO22X1 U171 ( .IN1(neighborCount[3]), .IN2(n84), .IN3(n85), .IN4(data_in[3]), 
        .Q(n181) );
  AO22X1 U172 ( .IN1(neighborCount[2]), .IN2(n84), .IN3(n85), .IN4(data_in[2]), 
        .Q(n182) );
  AO22X1 U173 ( .IN1(neighborCount[1]), .IN2(n84), .IN3(n85), .IN4(data_in[1]), 
        .Q(n183) );
  AO22X1 U174 ( .IN1(neighborCount[0]), .IN2(n84), .IN3(n85), .IN4(data_in[0]), 
        .Q(n184) );
  AO22X1 U175 ( .IN1(neighborID[15]), .IN2(n87), .IN3(n53), .IN4(data_in[15]), 
        .Q(n185) );
  AO22X1 U176 ( .IN1(neighborID[14]), .IN2(n87), .IN3(n53), .IN4(data_in[14]), 
        .Q(n186) );
  AO22X1 U177 ( .IN1(neighborID[13]), .IN2(n87), .IN3(n53), .IN4(data_in[13]), 
        .Q(n187) );
  AO22X1 U178 ( .IN1(neighborID[12]), .IN2(n87), .IN3(n53), .IN4(data_in[12]), 
        .Q(n188) );
  AO22X1 U179 ( .IN1(neighborID[11]), .IN2(n87), .IN3(n53), .IN4(data_in[11]), 
        .Q(n189) );
  AO22X1 U180 ( .IN1(neighborID[10]), .IN2(n87), .IN3(n53), .IN4(data_in[10]), 
        .Q(n190) );
  AO22X1 U181 ( .IN1(neighborID[9]), .IN2(n87), .IN3(n53), .IN4(data_in[9]), 
        .Q(n191) );
  AO22X1 U182 ( .IN1(neighborID[8]), .IN2(n87), .IN3(n53), .IN4(data_in[8]), 
        .Q(n192) );
  AO22X1 U183 ( .IN1(neighborID[7]), .IN2(n87), .IN3(n53), .IN4(data_in[7]), 
        .Q(n193) );
  AO22X1 U184 ( .IN1(neighborID[6]), .IN2(n87), .IN3(n53), .IN4(data_in[6]), 
        .Q(n194) );
  AO22X1 U185 ( .IN1(neighborID[5]), .IN2(n87), .IN3(n53), .IN4(data_in[5]), 
        .Q(n195) );
  AO22X1 U186 ( .IN1(neighborID[4]), .IN2(n87), .IN3(n53), .IN4(data_in[4]), 
        .Q(n196) );
  AO22X1 U187 ( .IN1(neighborID[3]), .IN2(n87), .IN3(n53), .IN4(data_in[3]), 
        .Q(n197) );
  AO22X1 U188 ( .IN1(neighborID[2]), .IN2(n87), .IN3(n53), .IN4(data_in[2]), 
        .Q(n198) );
  AO22X1 U189 ( .IN1(neighborID[1]), .IN2(n87), .IN3(n53), .IN4(data_in[1]), 
        .Q(n199) );
  AO22X1 U190 ( .IN1(clusterID[15]), .IN2(n88), .IN3(n54), .IN4(data_in[15]), 
        .Q(n200) );
  AO22X1 U191 ( .IN1(clusterID[14]), .IN2(n88), .IN3(n54), .IN4(data_in[14]), 
        .Q(n201) );
  AO22X1 U192 ( .IN1(clusterID[13]), .IN2(n88), .IN3(n54), .IN4(data_in[13]), 
        .Q(n202) );
  AO22X1 U193 ( .IN1(clusterID[12]), .IN2(n88), .IN3(n54), .IN4(data_in[12]), 
        .Q(n203) );
  AO22X1 U194 ( .IN1(clusterID[11]), .IN2(n88), .IN3(n54), .IN4(data_in[11]), 
        .Q(n204) );
  AO22X1 U195 ( .IN1(clusterID[10]), .IN2(n88), .IN3(n54), .IN4(data_in[10]), 
        .Q(n205) );
  AO22X1 U196 ( .IN1(clusterID[9]), .IN2(n88), .IN3(n54), .IN4(data_in[9]), 
        .Q(n206) );
  AO22X1 U197 ( .IN1(clusterID[8]), .IN2(n88), .IN3(n54), .IN4(data_in[8]), 
        .Q(n207) );
  AO22X1 U198 ( .IN1(clusterID[7]), .IN2(n88), .IN3(n54), .IN4(data_in[7]), 
        .Q(n208) );
  AO22X1 U199 ( .IN1(clusterID[6]), .IN2(n88), .IN3(n54), .IN4(data_in[6]), 
        .Q(n209) );
  AO22X1 U200 ( .IN1(clusterID[5]), .IN2(n88), .IN3(n54), .IN4(data_in[5]), 
        .Q(n210) );
  AO22X1 U201 ( .IN1(clusterID[4]), .IN2(n88), .IN3(n54), .IN4(data_in[4]), 
        .Q(n211) );
  AO22X1 U202 ( .IN1(clusterID[3]), .IN2(n88), .IN3(n54), .IN4(data_in[3]), 
        .Q(n212) );
  AO22X1 U203 ( .IN1(clusterID[2]), .IN2(n88), .IN3(n54), .IN4(data_in[2]), 
        .Q(n213) );
  AO22X1 U204 ( .IN1(clusterID[1]), .IN2(n88), .IN3(n54), .IN4(data_in[1]), 
        .Q(n214) );
  AO22X1 U205 ( .IN1(clusterID[0]), .IN2(n88), .IN3(n54), .IN4(data_in[0]), 
        .Q(n215) );
  AO221X1 U206 ( .IN1(n90), .IN2(n91), .IN3(nrst), .IN4(n92), .IN5(n93), .Q(
        n216) );
  NAND3X0 U207 ( .IN1(n77), .IN2(n38), .IN3(n89), .QN(n92) );
  OR2X1 U208 ( .IN1(N204), .IN2(n332), .Q(n91) );
  AO21X1 U209 ( .IN1(nrst), .IN2(n95), .IN3(n90), .Q(n217) );
  AO221X1 U210 ( .IN1(nrst), .IN2(n96), .IN3(n90), .IN4(n94), .IN5(n93), .Q(
        n218) );
  AND4X1 U211 ( .IN1(n39), .IN2(n223), .IN3(n97), .IN4(n98), .Q(n93) );
  NOR4X0 U212 ( .IN1(n69), .IN2(n334), .IN3(n333), .IN4(n95), .QN(n98) );
  NAND3X0 U213 ( .IN1(n76), .IN2(n38), .IN3(n86), .QN(n95) );
  NAND3X0 U214 ( .IN1(n30), .IN2(n29), .IN3(n99), .QN(n76) );
  NAND3X0 U215 ( .IN1(n101), .IN2(state[2]), .IN3(state[1]), .QN(n38) );
  AND3X1 U216 ( .IN1(n86), .IN2(n89), .IN3(n102), .Q(n75) );
  NAND3X0 U217 ( .IN1(state[2]), .IN2(n30), .IN3(n101), .QN(n89) );
  NAND3X0 U218 ( .IN1(n101), .IN2(n29), .IN3(state[1]), .QN(n86) );
  NAND4X0 U219 ( .IN1(nrst), .IN2(n104), .IN3(n105), .IN4(n100), .QN(n219) );
  NAND3X0 U220 ( .IN1(state[2]), .IN2(n99), .IN3(state[1]), .QN(n100) );
  AO22X1 U221 ( .IN1(neighborID[0]), .IN2(n87), .IN3(n53), .IN4(data_in[0]), 
        .Q(n220) );
  NAND3X0 U222 ( .IN1(n99), .IN2(n29), .IN3(state[1]), .QN(n77) );
  AO21X1 U223 ( .IN1(en), .IN2(n41), .IN3(n328), .Q(n81) );
  NAND3X0 U224 ( .IN1(n30), .IN2(n29), .IN3(n31), .QN(n103) );
  NAND3X0 U225 ( .IN1(n99), .IN2(n30), .IN3(state[2]), .QN(n68) );
  AO22X1 U226 ( .IN1(N151), .IN2(n222), .IN3(N80), .IN4(n223), .Q(N203) );
  AO22X1 U227 ( .IN1(N152), .IN2(n222), .IN3(N81), .IN4(n223), .Q(N202) );
  AO22X1 U228 ( .IN1(N136), .IN2(n222), .IN3(i[2]), .IN4(n223), .Q(N201) );
  AO22X1 U229 ( .IN1(N137), .IN2(n222), .IN3(i[3]), .IN4(n223), .Q(N200) );
  AO22X1 U230 ( .IN1(N138), .IN2(n222), .IN3(i[4]), .IN4(n223), .Q(N199) );
  AO22X1 U231 ( .IN1(N139), .IN2(n222), .IN3(i[5]), .IN4(n223), .Q(N198) );
  AO22X1 U232 ( .IN1(N140), .IN2(n222), .IN3(i[6]), .IN4(n223), .Q(N197) );
  AO22X1 U233 ( .IN1(N141), .IN2(n222), .IN3(i[7]), .IN4(n223), .Q(N196) );
  AO22X1 U234 ( .IN1(N142), .IN2(n222), .IN3(i[8]), .IN4(n223), .Q(N195) );
  AO22X1 U235 ( .IN1(N143), .IN2(n222), .IN3(i[9]), .IN4(n223), .Q(N194) );
  AO22X1 U236 ( .IN1(N144), .IN2(n222), .IN3(i[10]), .IN4(n223), .Q(N193) );
  AO22X1 U237 ( .IN1(N145), .IN2(n222), .IN3(i[11]), .IN4(n223), .Q(N192) );
  AO22X1 U238 ( .IN1(N146), .IN2(n222), .IN3(i[12]), .IN4(n223), .Q(N191) );
  AO22X1 U239 ( .IN1(N147), .IN2(n222), .IN3(i[13]), .IN4(n223), .Q(N190) );
  AO22X1 U240 ( .IN1(N148), .IN2(n222), .IN3(i[14]), .IN4(n223), .Q(N189) );
  AO22X1 U241 ( .IN1(N149), .IN2(n222), .IN3(i[15]), .IN4(n223), .Q(N188) );
  neighborSinkInOtherCluster_DW01_inc_0 add_90 ( .A({i[15:2], N81, N80}), 
        .SUM({N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N152, N151}) );
  neighborSinkInOtherCluster_DW01_inc_1 add_85 ( .A({j[15:2], N92, N91}), 
        .SUM({N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, 
        N109, N108, N107, N123, N122}) );
  DFFX1 done_buf_reg ( .D(n107), .CLK(clock), .Q(done) );
  DFFX1 \knownSinkCount_reg[15]  ( .D(n153), .CLK(clock), .Q(
        knownSinkCount[15]) );
  DFFX1 \knownSinkCount_reg[14]  ( .D(n154), .CLK(clock), .Q(
        knownSinkCount[14]) );
  DFFX1 \knownSinkCount_reg[13]  ( .D(n155), .CLK(clock), .Q(
        knownSinkCount[13]) );
  DFFX1 \knownSinkCount_reg[12]  ( .D(n156), .CLK(clock), .Q(
        knownSinkCount[12]) );
  DFFX1 \knownSinkCount_reg[11]  ( .D(n157), .CLK(clock), .Q(
        knownSinkCount[11]) );
  DFFX1 \knownSinkCount_reg[10]  ( .D(n158), .CLK(clock), .Q(
        knownSinkCount[10]) );
  DFFX1 \knownSinkCount_reg[9]  ( .D(n159), .CLK(clock), .Q(knownSinkCount[9])
         );
  DFFX1 \knownSinkCount_reg[8]  ( .D(n160), .CLK(clock), .Q(knownSinkCount[8])
         );
  DFFX1 \knownSinkCount_reg[7]  ( .D(n161), .CLK(clock), .Q(knownSinkCount[7])
         );
  DFFX1 \knownSinkCount_reg[6]  ( .D(n162), .CLK(clock), .Q(knownSinkCount[6])
         );
  DFFX1 \knownSinkCount_reg[5]  ( .D(n163), .CLK(clock), .Q(knownSinkCount[5])
         );
  DFFX1 \knownSinkCount_reg[4]  ( .D(n164), .CLK(clock), .Q(knownSinkCount[4])
         );
  DFFX1 \knownSinkCount_reg[3]  ( .D(n165), .CLK(clock), .Q(knownSinkCount[3])
         );
  DFFX1 \knownSinkCount_reg[2]  ( .D(n166), .CLK(clock), .Q(knownSinkCount[2])
         );
  DFFX1 \knownSinkCount_reg[1]  ( .D(n167), .CLK(clock), .Q(knownSinkCount[1]), 
        .QN(n298) );
  DFFX1 \knownSinkCount_reg[0]  ( .D(n168), .CLK(clock), .Q(knownSinkCount[0]), 
        .QN(n297) );
  DFFX1 \neighborCount_reg[15]  ( .D(n169), .CLK(clock), .Q(neighborCount[15])
         );
  DFFX1 \neighborCount_reg[14]  ( .D(n170), .CLK(clock), .Q(neighborCount[14])
         );
  DFFX1 \neighborCount_reg[13]  ( .D(n171), .CLK(clock), .Q(neighborCount[13])
         );
  DFFX1 \neighborCount_reg[12]  ( .D(n172), .CLK(clock), .Q(neighborCount[12])
         );
  DFFX1 \neighborCount_reg[11]  ( .D(n173), .CLK(clock), .Q(neighborCount[11])
         );
  DFFX1 \neighborCount_reg[10]  ( .D(n174), .CLK(clock), .Q(neighborCount[10])
         );
  DFFX1 \neighborCount_reg[9]  ( .D(n175), .CLK(clock), .Q(neighborCount[9])
         );
  DFFX1 \neighborCount_reg[8]  ( .D(n176), .CLK(clock), .Q(neighborCount[8])
         );
  DFFX1 \neighborCount_reg[7]  ( .D(n177), .CLK(clock), .Q(neighborCount[7])
         );
  DFFX1 \neighborCount_reg[6]  ( .D(n178), .CLK(clock), .Q(neighborCount[6])
         );
  DFFX1 \neighborCount_reg[5]  ( .D(n179), .CLK(clock), .Q(neighborCount[5])
         );
  DFFX1 \neighborCount_reg[4]  ( .D(n180), .CLK(clock), .Q(neighborCount[4])
         );
  DFFX1 \neighborCount_reg[3]  ( .D(n181), .CLK(clock), .Q(neighborCount[3])
         );
  DFFX1 \neighborCount_reg[2]  ( .D(n182), .CLK(clock), .Q(neighborCount[2])
         );
  DFFX1 \neighborCount_reg[1]  ( .D(n183), .CLK(clock), .Q(neighborCount[1]), 
        .QN(n322) );
  DFFX1 \neighborCount_reg[0]  ( .D(n184), .CLK(clock), .Q(neighborCount[0]), 
        .QN(n323) );
  DFFX1 \clusterID_reg[15]  ( .D(n200), .CLK(clock), .Q(clusterID[15]) );
  DFFX1 \clusterID_reg[14]  ( .D(n201), .CLK(clock), .Q(clusterID[14]) );
  DFFX1 \clusterID_reg[13]  ( .D(n202), .CLK(clock), .Q(clusterID[13]) );
  DFFX1 \clusterID_reg[12]  ( .D(n203), .CLK(clock), .Q(clusterID[12]) );
  DFFX1 \clusterID_reg[11]  ( .D(n204), .CLK(clock), .Q(clusterID[11]) );
  DFFX1 \clusterID_reg[10]  ( .D(n205), .CLK(clock), .Q(clusterID[10]) );
  DFFX1 \clusterID_reg[9]  ( .D(n206), .CLK(clock), .Q(clusterID[9]) );
  DFFX1 \clusterID_reg[8]  ( .D(n207), .CLK(clock), .Q(clusterID[8]) );
  DFFX1 \clusterID_reg[7]  ( .D(n208), .CLK(clock), .Q(clusterID[7]) );
  DFFX1 \clusterID_reg[6]  ( .D(n209), .CLK(clock), .Q(clusterID[6]) );
  DFFX1 \clusterID_reg[5]  ( .D(n210), .CLK(clock), .Q(clusterID[5]) );
  DFFX1 \clusterID_reg[4]  ( .D(n211), .CLK(clock), .Q(clusterID[4]) );
  DFFX1 \clusterID_reg[3]  ( .D(n212), .CLK(clock), .Q(clusterID[3]) );
  DFFX1 \clusterID_reg[2]  ( .D(n213), .CLK(clock), .Q(clusterID[2]) );
  DFFX1 \clusterID_reg[1]  ( .D(n214), .CLK(clock), .Q(clusterID[1]), .QN(n272) );
  DFFX1 \clusterID_reg[0]  ( .D(n215), .CLK(clock), .Q(clusterID[0]), .QN(n271) );
  DFFX1 \neighborID_reg[15]  ( .D(n185), .CLK(clock), .Q(neighborID[15]) );
  DFFX1 \neighborID_reg[14]  ( .D(n186), .CLK(clock), .Q(neighborID[14]) );
  DFFX1 \neighborID_reg[13]  ( .D(n187), .CLK(clock), .Q(neighborID[13]) );
  DFFX1 \neighborID_reg[12]  ( .D(n188), .CLK(clock), .Q(neighborID[12]) );
  DFFX1 \neighborID_reg[11]  ( .D(n189), .CLK(clock), .Q(neighborID[11]) );
  DFFX1 \neighborID_reg[10]  ( .D(n190), .CLK(clock), .Q(neighborID[10]) );
  DFFX1 \neighborID_reg[9]  ( .D(n191), .CLK(clock), .Q(neighborID[9]) );
  DFFX1 \neighborID_reg[8]  ( .D(n192), .CLK(clock), .Q(neighborID[8]) );
  DFFX1 \neighborID_reg[7]  ( .D(n193), .CLK(clock), .Q(neighborID[7]) );
  DFFX1 \neighborID_reg[6]  ( .D(n194), .CLK(clock), .Q(neighborID[6]) );
  DFFX1 \neighborID_reg[5]  ( .D(n195), .CLK(clock), .Q(neighborID[5]) );
  DFFX1 \neighborID_reg[4]  ( .D(n196), .CLK(clock), .Q(neighborID[4]) );
  DFFX1 \neighborID_reg[3]  ( .D(n197), .CLK(clock), .Q(neighborID[3]) );
  DFFX1 \neighborID_reg[2]  ( .D(n198), .CLK(clock), .Q(neighborID[2]) );
  DFFX1 \neighborID_reg[1]  ( .D(n199), .CLK(clock), .Q(neighborID[1]), .QN(
        n246) );
  DFFX1 \neighborID_reg[0]  ( .D(n220), .CLK(clock), .Q(neighborID[0]) );
  DFFX1 \j_reg[15]  ( .D(n137), .CLK(clock), .Q(j[15]) );
  DFFX1 \j_reg[14]  ( .D(n138), .CLK(clock), .Q(j[14]) );
  DFFX1 \j_reg[13]  ( .D(n139), .CLK(clock), .Q(j[13]) );
  DFFX1 \j_reg[12]  ( .D(n140), .CLK(clock), .Q(j[12]) );
  DFFX1 \j_reg[11]  ( .D(n141), .CLK(clock), .Q(j[11]) );
  DFFX1 \j_reg[10]  ( .D(n142), .CLK(clock), .Q(j[10]) );
  DFFX1 \j_reg[9]  ( .D(n143), .CLK(clock), .Q(j[9]) );
  DFFX1 \j_reg[8]  ( .D(n144), .CLK(clock), .Q(j[8]) );
  DFFX1 \j_reg[7]  ( .D(n145), .CLK(clock), .Q(j[7]) );
  DFFX1 \j_reg[6]  ( .D(n146), .CLK(clock), .Q(j[6]) );
  DFFX1 \j_reg[5]  ( .D(n147), .CLK(clock), .Q(j[5]) );
  DFFX1 \j_reg[4]  ( .D(n148), .CLK(clock), .Q(j[4]) );
  DFFX1 \j_reg[3]  ( .D(n149), .CLK(clock), .Q(j[3]) );
  DFFX1 \j_reg[2]  ( .D(n150), .CLK(clock), .Q(j[2]), .QN(N93) );
  DFFX1 \j_reg[1]  ( .D(n151), .CLK(clock), .Q(N92) );
  DFFX1 \j_reg[0]  ( .D(n152), .CLK(clock), .Q(N91) );
  DFFX1 forAggregation_buf_reg ( .D(n108), .CLK(clock), .Q(forAggregation) );
  DFFX1 \address_count_reg[0]  ( .D(n221), .CLK(clock), .Q(address[0]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n120), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \i_reg[15]  ( .D(n136), .CLK(clock), .Q(i[15]) );
  DFFX1 \i_reg[14]  ( .D(n121), .CLK(clock), .Q(i[14]) );
  DFFX1 \i_reg[13]  ( .D(n122), .CLK(clock), .Q(i[13]) );
  DFFX1 \i_reg[12]  ( .D(n123), .CLK(clock), .Q(i[12]) );
  DFFX1 \i_reg[11]  ( .D(n124), .CLK(clock), .Q(i[11]) );
  DFFX1 \i_reg[10]  ( .D(n125), .CLK(clock), .Q(i[10]) );
  DFFX1 \i_reg[9]  ( .D(n126), .CLK(clock), .Q(i[9]) );
  DFFX1 \i_reg[8]  ( .D(n127), .CLK(clock), .Q(i[8]) );
  DFFX1 \i_reg[7]  ( .D(n128), .CLK(clock), .Q(i[7]) );
  DFFX1 \i_reg[6]  ( .D(n129), .CLK(clock), .Q(i[6]) );
  DFFX1 \i_reg[5]  ( .D(n130), .CLK(clock), .Q(i[5]) );
  DFFX1 \i_reg[4]  ( .D(n131), .CLK(clock), .Q(i[4]) );
  DFFX1 \i_reg[3]  ( .D(n132), .CLK(clock), .Q(i[3]) );
  DFFX1 \i_reg[2]  ( .D(n133), .CLK(clock), .Q(i[2]), .QN(N82) );
  DFFX1 \i_reg[1]  ( .D(n134), .CLK(clock), .Q(N81) );
  DFFX1 \i_reg[0]  ( .D(n135), .CLK(clock), .Q(N80) );
  DFFX1 \address_count_reg[1]  ( .D(n118), .CLK(clock), .Q(address[1]) );
  DFFX1 wr_en_buf_reg ( .D(n106), .CLK(clock), .Q(wr_en) );
  DFFX1 \address_count_reg[2]  ( .D(n117), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[8]  ( .D(n111), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[5]  ( .D(n114), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n115), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[10]  ( .D(n109), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n110), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[7]  ( .D(n112), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[6]  ( .D(n113), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[3]  ( .D(n116), .CLK(clock), .Q(address[3]) );
  NOR2X0 U242 ( .IN1(n327), .IN2(n332), .QN(n74) );
  INVX0 U243 ( .INP(n36), .ZN(n327) );
  NOR2X0 U244 ( .IN1(n327), .IN2(n222), .QN(n80) );
  NOR2X0 U245 ( .IN1(n327), .IN2(n78), .QN(n79) );
  INVX0 U246 ( .INP(n43), .ZN(n324) );
  INVX0 U247 ( .INP(n94), .ZN(n332) );
  INVX0 U248 ( .INP(n59), .ZN(n326) );
  INVX0 U249 ( .INP(n222), .ZN(n223) );
  NOR2X0 U250 ( .IN1(n89), .IN2(n328), .QN(n54) );
  NOR2X0 U251 ( .IN1(n77), .IN2(n328), .QN(n53) );
  NOR2X0 U252 ( .IN1(n76), .IN2(n328), .QN(n83) );
  NOR2X0 U253 ( .IN1(n86), .IN2(n328), .QN(n85) );
  NOR2X0 U254 ( .IN1(n81), .IN2(n335), .QN(n82) );
  NOR2X0 U255 ( .IN1(n81), .IN2(n337), .QN(n88) );
  NOR2X0 U256 ( .IN1(n81), .IN2(n336), .QN(n84) );
  NOR2X0 U257 ( .IN1(n81), .IN2(n333), .QN(n87) );
  OA21X1 U258 ( .IN1(n223), .IN2(n68), .IN3(n325), .Q(n78) );
  NOR2X0 U259 ( .IN1(n328), .IN2(n68), .QN(n36) );
  AND2X1 U260 ( .IN1(n325), .IN2(n68), .Q(n42) );
  NOR2X0 U261 ( .IN1(n68), .IN2(n332), .QN(n45) );
  INVX0 U262 ( .INP(n81), .ZN(n325) );
  NOR2X0 U263 ( .IN1(n327), .IN2(n93), .QN(n90) );
  NAND2X1 U264 ( .IN1(N103), .IN2(N102), .QN(n94) );
  NBUFFX2 U265 ( .INP(N132), .Z(n222) );
  INVX0 U266 ( .INP(N107), .ZN(N124) );
  INVX0 U267 ( .INP(N136), .ZN(N153) );
  INVX0 U268 ( .INP(N202), .ZN(n321) );
  INVX0 U269 ( .INP(N123), .ZN(n296) );
  INVX0 U270 ( .INP(n77), .ZN(n333) );
  INVX0 U271 ( .INP(n89), .ZN(n337) );
  INVX0 U272 ( .INP(n76), .ZN(n335) );
  INVX0 U273 ( .INP(n86), .ZN(n336) );
  INVX0 U274 ( .INP(n100), .ZN(n334) );
  INVX0 U275 ( .INP(nrst), .ZN(n328) );
  NOR2X0 U276 ( .IN1(state[3]), .IN2(N204), .QN(n97) );
  NAND2X1 U277 ( .IN1(start), .IN2(n69), .QN(n102) );
  OA21X1 U278 ( .IN1(n94), .IN2(n68), .IN3(nrst), .Q(n39) );
  NAND2X1 U279 ( .IN1(n75), .IN2(n38), .QN(n96) );
  AND2X1 U280 ( .IN1(address[0]), .IN2(n324), .Q(n221) );
  INVX0 U281 ( .INP(data_in[1]), .ZN(n248) );
  INVX0 U282 ( .INP(n37), .ZN(n330) );
  NAND2X1 U283 ( .IN1(en), .IN2(n41), .QN(n40) );
  NAND2X1 U284 ( .IN1(N82), .IN2(n333), .QN(n65) );
  INVX0 U285 ( .INP(n39), .ZN(n329) );
  NAND2X1 U286 ( .IN1(state[3]), .IN2(n103), .QN(n104) );
  NAND2X1 U287 ( .IN1(n41), .IN2(n331), .QN(n105) );
  INVX0 U288 ( .INP(en), .ZN(n331) );
  INVX0 U289 ( .INP(data_in[0]), .ZN(n247) );
  INVX0 U290 ( .INP(MY_CLUSTER_ID[1]), .ZN(n273) );
  NOR2X0 U291 ( .IN1(n23), .IN2(n103), .QN(n41) );
  NOR2X0 U292 ( .IN1(n103), .IN2(state[3]), .QN(n69) );
  NOR2X0 U293 ( .IN1(n31), .IN2(state[3]), .QN(n99) );
  NOR2X0 U294 ( .IN1(state[3]), .IN2(state[0]), .QN(n101) );
  XOR2X1 U295 ( .IN1(i[9]), .IN2(\add_66/carry[10] ), .Q(N89) );
  XOR2X1 U296 ( .IN1(j[9]), .IN2(\add_72/carry[10] ), .Q(N100) );
  XOR2X1 U297 ( .IN1(N114), .IN2(\add_86/carry[10] ), .Q(N131) );
  XOR2X1 U298 ( .IN1(N143), .IN2(\add_92/carry[10] ), .Q(N160) );
  AND2X1 U299 ( .IN1(\add_66/carry[9] ), .IN2(i[8]), .Q(\add_66/carry[10] ) );
  XOR2X1 U300 ( .IN1(i[8]), .IN2(\add_66/carry[9] ), .Q(N88) );
  AND2X1 U301 ( .IN1(\add_72/carry[9] ), .IN2(j[8]), .Q(\add_72/carry[10] ) );
  XOR2X1 U302 ( .IN1(j[8]), .IN2(\add_72/carry[9] ), .Q(N99) );
  AND2X1 U303 ( .IN1(\add_86/carry[9] ), .IN2(N113), .Q(\add_86/carry[10] ) );
  XOR2X1 U304 ( .IN1(N113), .IN2(\add_86/carry[9] ), .Q(N130) );
  AND2X1 U305 ( .IN1(\add_92/carry[9] ), .IN2(N142), .Q(\add_92/carry[10] ) );
  XOR2X1 U306 ( .IN1(N142), .IN2(\add_92/carry[9] ), .Q(N159) );
  AND2X1 U307 ( .IN1(\add_86/carry[8] ), .IN2(N112), .Q(\add_86/carry[9] ) );
  XOR2X1 U308 ( .IN1(N112), .IN2(\add_86/carry[8] ), .Q(N129) );
  AND2X1 U309 ( .IN1(\add_72/carry[8] ), .IN2(j[7]), .Q(\add_72/carry[9] ) );
  XOR2X1 U310 ( .IN1(j[7]), .IN2(\add_72/carry[8] ), .Q(N98) );
  AND2X1 U311 ( .IN1(\add_66/carry[8] ), .IN2(i[7]), .Q(\add_66/carry[9] ) );
  XOR2X1 U312 ( .IN1(i[7]), .IN2(\add_66/carry[8] ), .Q(N87) );
  AND2X1 U313 ( .IN1(\add_92/carry[8] ), .IN2(N141), .Q(\add_92/carry[9] ) );
  XOR2X1 U314 ( .IN1(N141), .IN2(\add_92/carry[8] ), .Q(N158) );
  OR2X1 U315 ( .IN1(i[6]), .IN2(\add_66/carry[7] ), .Q(\add_66/carry[8] ) );
  XNOR2X1 U316 ( .IN1(\add_66/carry[7] ), .IN2(i[6]), .Q(N86) );
  AND2X1 U317 ( .IN1(\add_72/carry[7] ), .IN2(j[6]), .Q(\add_72/carry[8] ) );
  XOR2X1 U318 ( .IN1(j[6]), .IN2(\add_72/carry[7] ), .Q(N97) );
  AND2X1 U319 ( .IN1(\add_86/carry[7] ), .IN2(N111), .Q(\add_86/carry[8] ) );
  XOR2X1 U320 ( .IN1(N111), .IN2(\add_86/carry[7] ), .Q(N128) );
  AND2X1 U321 ( .IN1(\add_92/carry[7] ), .IN2(N140), .Q(\add_92/carry[8] ) );
  XOR2X1 U322 ( .IN1(N140), .IN2(\add_92/carry[7] ), .Q(N157) );
  AND2X1 U323 ( .IN1(\add_86/carry[6] ), .IN2(N110), .Q(\add_86/carry[7] ) );
  XOR2X1 U324 ( .IN1(N110), .IN2(\add_86/carry[6] ), .Q(N127) );
  OR2X1 U325 ( .IN1(N139), .IN2(\add_92/carry[6] ), .Q(\add_92/carry[7] ) );
  XNOR2X1 U326 ( .IN1(\add_92/carry[6] ), .IN2(N139), .Q(N156) );
  OR2X1 U327 ( .IN1(i[5]), .IN2(\add_66/carry[6] ), .Q(\add_66/carry[7] ) );
  XNOR2X1 U328 ( .IN1(\add_66/carry[6] ), .IN2(i[5]), .Q(N85) );
  AND2X1 U329 ( .IN1(\add_72/carry[6] ), .IN2(j[5]), .Q(\add_72/carry[7] ) );
  XOR2X1 U330 ( .IN1(j[5]), .IN2(\add_72/carry[6] ), .Q(N96) );
  AND2X1 U331 ( .IN1(\add_86/carry[5] ), .IN2(N109), .Q(\add_86/carry[6] ) );
  XOR2X1 U332 ( .IN1(N109), .IN2(\add_86/carry[5] ), .Q(N126) );
  AND2X1 U333 ( .IN1(\add_72/carry[5] ), .IN2(j[4]), .Q(\add_72/carry[6] ) );
  XOR2X1 U334 ( .IN1(j[4]), .IN2(\add_72/carry[5] ), .Q(N95) );
  AND2X1 U335 ( .IN1(\add_66/carry[5] ), .IN2(i[4]), .Q(\add_66/carry[6] ) );
  XOR2X1 U336 ( .IN1(i[4]), .IN2(\add_66/carry[5] ), .Q(N84) );
  AND2X1 U337 ( .IN1(\add_92/carry[5] ), .IN2(N138), .Q(\add_92/carry[6] ) );
  XOR2X1 U338 ( .IN1(N138), .IN2(\add_92/carry[5] ), .Q(N155) );
  AND2X1 U339 ( .IN1(N107), .IN2(N108), .Q(\add_86/carry[5] ) );
  XOR2X1 U340 ( .IN1(N108), .IN2(N107), .Q(N125) );
  AND2X1 U341 ( .IN1(j[2]), .IN2(j[3]), .Q(\add_72/carry[5] ) );
  XOR2X1 U342 ( .IN1(j[3]), .IN2(j[2]), .Q(N94) );
  AND2X1 U343 ( .IN1(i[2]), .IN2(i[3]), .Q(\add_66/carry[5] ) );
  XOR2X1 U344 ( .IN1(i[3]), .IN2(i[2]), .Q(N83) );
  AND2X1 U345 ( .IN1(N136), .IN2(N137), .Q(\add_92/carry[5] ) );
  XOR2X1 U346 ( .IN1(N137), .IN2(N136), .Q(N154) );
  XOR2X1 U347 ( .IN1(data_in[15]), .IN2(neighborID[15]), .Q(n229) );
  XOR2X1 U348 ( .IN1(data_in[2]), .IN2(neighborID[2]), .Q(n228) );
  NOR2X0 U349 ( .IN1(n247), .IN2(neighborID[0]), .QN(n224) );
  OA22X1 U350 ( .IN1(data_in[1]), .IN2(n224), .IN3(n224), .IN4(n246), .Q(n227)
         );
  AND2X1 U351 ( .IN1(neighborID[0]), .IN2(n247), .Q(n225) );
  OA22X1 U352 ( .IN1(n225), .IN2(n248), .IN3(neighborID[1]), .IN4(n225), .Q(
        n226) );
  OR4X1 U353 ( .IN1(n229), .IN2(n228), .IN3(n227), .IN4(n226), .Q(n245) );
  XNOR2X1 U354 ( .IN1(data_in[6]), .IN2(neighborID[6]), .Q(n233) );
  XNOR2X1 U355 ( .IN1(data_in[5]), .IN2(neighborID[5]), .Q(n232) );
  XNOR2X1 U356 ( .IN1(data_in[4]), .IN2(neighborID[4]), .Q(n231) );
  XNOR2X1 U357 ( .IN1(data_in[3]), .IN2(neighborID[3]), .Q(n230) );
  NAND4X0 U358 ( .IN1(n233), .IN2(n232), .IN3(n231), .IN4(n230), .QN(n244) );
  XNOR2X1 U359 ( .IN1(data_in[10]), .IN2(neighborID[10]), .Q(n237) );
  XNOR2X1 U360 ( .IN1(data_in[9]), .IN2(neighborID[9]), .Q(n236) );
  XNOR2X1 U361 ( .IN1(data_in[8]), .IN2(neighborID[8]), .Q(n235) );
  XNOR2X1 U362 ( .IN1(data_in[7]), .IN2(neighborID[7]), .Q(n234) );
  NAND4X0 U363 ( .IN1(n237), .IN2(n236), .IN3(n235), .IN4(n234), .QN(n243) );
  XNOR2X1 U364 ( .IN1(data_in[14]), .IN2(neighborID[14]), .Q(n241) );
  XNOR2X1 U365 ( .IN1(data_in[13]), .IN2(neighborID[13]), .Q(n240) );
  XNOR2X1 U366 ( .IN1(data_in[12]), .IN2(neighborID[12]), .Q(n239) );
  XNOR2X1 U367 ( .IN1(data_in[11]), .IN2(neighborID[11]), .Q(n238) );
  NAND4X0 U368 ( .IN1(n241), .IN2(n240), .IN3(n239), .IN4(n238), .QN(n242) );
  NOR4X0 U369 ( .IN1(n245), .IN2(n244), .IN3(n243), .IN4(n242), .QN(N102) );
  XOR2X1 U370 ( .IN1(MY_CLUSTER_ID[12]), .IN2(clusterID[12]), .Q(n252) );
  XOR2X1 U371 ( .IN1(MY_CLUSTER_ID[13]), .IN2(clusterID[13]), .Q(n251) );
  XOR2X1 U372 ( .IN1(MY_CLUSTER_ID[14]), .IN2(clusterID[14]), .Q(n250) );
  XOR2X1 U373 ( .IN1(MY_CLUSTER_ID[15]), .IN2(clusterID[15]), .Q(n249) );
  NOR4X0 U374 ( .IN1(n252), .IN2(n251), .IN3(n250), .IN4(n249), .QN(n270) );
  XOR2X1 U375 ( .IN1(MY_CLUSTER_ID[8]), .IN2(clusterID[8]), .Q(n256) );
  XOR2X1 U376 ( .IN1(MY_CLUSTER_ID[9]), .IN2(clusterID[9]), .Q(n255) );
  XOR2X1 U377 ( .IN1(MY_CLUSTER_ID[10]), .IN2(clusterID[10]), .Q(n254) );
  XOR2X1 U378 ( .IN1(MY_CLUSTER_ID[11]), .IN2(clusterID[11]), .Q(n253) );
  NOR4X0 U379 ( .IN1(n256), .IN2(n255), .IN3(n254), .IN4(n253), .QN(n269) );
  XOR2X1 U380 ( .IN1(MY_CLUSTER_ID[4]), .IN2(clusterID[4]), .Q(n260) );
  XOR2X1 U381 ( .IN1(MY_CLUSTER_ID[5]), .IN2(clusterID[5]), .Q(n259) );
  XOR2X1 U382 ( .IN1(MY_CLUSTER_ID[6]), .IN2(clusterID[6]), .Q(n258) );
  XOR2X1 U383 ( .IN1(MY_CLUSTER_ID[7]), .IN2(clusterID[7]), .Q(n257) );
  NOR4X0 U384 ( .IN1(n260), .IN2(n259), .IN3(n258), .IN4(n257), .QN(n268) );
  NOR2X0 U385 ( .IN1(n271), .IN2(MY_CLUSTER_ID[0]), .QN(n261) );
  OA22X1 U386 ( .IN1(n261), .IN2(n273), .IN3(clusterID[1]), .IN4(n261), .Q(
        n266) );
  AND2X1 U387 ( .IN1(MY_CLUSTER_ID[0]), .IN2(n271), .Q(n262) );
  OA22X1 U388 ( .IN1(MY_CLUSTER_ID[1]), .IN2(n262), .IN3(n262), .IN4(n272), 
        .Q(n265) );
  XOR2X1 U389 ( .IN1(MY_CLUSTER_ID[2]), .IN2(clusterID[2]), .Q(n264) );
  XOR2X1 U390 ( .IN1(MY_CLUSTER_ID[3]), .IN2(clusterID[3]), .Q(n263) );
  NOR4X0 U391 ( .IN1(n266), .IN2(n265), .IN3(n264), .IN4(n263), .QN(n267) );
  NAND4X0 U392 ( .IN1(n270), .IN2(n269), .IN3(n268), .IN4(n267), .QN(N103) );
  XOR2X1 U393 ( .IN1(knownSinkCount[15]), .IN2(N120), .Q(n279) );
  XOR2X1 U394 ( .IN1(knownSinkCount[2]), .IN2(N107), .Q(n278) );
  NOR2X0 U395 ( .IN1(n297), .IN2(N122), .QN(n274) );
  OA22X1 U396 ( .IN1(knownSinkCount[1]), .IN2(n274), .IN3(n274), .IN4(n296), 
        .Q(n277) );
  AND2X1 U397 ( .IN1(N122), .IN2(n297), .Q(n275) );
  OA22X1 U398 ( .IN1(n275), .IN2(n298), .IN3(N123), .IN4(n275), .Q(n276) );
  OR4X1 U399 ( .IN1(n279), .IN2(n278), .IN3(n277), .IN4(n276), .Q(n295) );
  XNOR2X1 U400 ( .IN1(knownSinkCount[6]), .IN2(N111), .Q(n283) );
  XNOR2X1 U401 ( .IN1(knownSinkCount[5]), .IN2(N110), .Q(n282) );
  XNOR2X1 U402 ( .IN1(knownSinkCount[4]), .IN2(N109), .Q(n281) );
  XNOR2X1 U403 ( .IN1(knownSinkCount[3]), .IN2(N108), .Q(n280) );
  NAND4X0 U404 ( .IN1(n283), .IN2(n282), .IN3(n281), .IN4(n280), .QN(n294) );
  XNOR2X1 U405 ( .IN1(knownSinkCount[10]), .IN2(N115), .Q(n287) );
  XNOR2X1 U406 ( .IN1(knownSinkCount[9]), .IN2(N114), .Q(n286) );
  XNOR2X1 U407 ( .IN1(knownSinkCount[8]), .IN2(N113), .Q(n285) );
  XNOR2X1 U408 ( .IN1(knownSinkCount[7]), .IN2(N112), .Q(n284) );
  NAND4X0 U409 ( .IN1(n287), .IN2(n286), .IN3(n285), .IN4(n284), .QN(n293) );
  XNOR2X1 U410 ( .IN1(knownSinkCount[14]), .IN2(N119), .Q(n291) );
  XNOR2X1 U411 ( .IN1(knownSinkCount[13]), .IN2(N118), .Q(n290) );
  XNOR2X1 U412 ( .IN1(knownSinkCount[12]), .IN2(N117), .Q(n289) );
  XNOR2X1 U413 ( .IN1(knownSinkCount[11]), .IN2(N116), .Q(n288) );
  NAND4X0 U414 ( .IN1(n291), .IN2(n290), .IN3(n289), .IN4(n288), .QN(n292) );
  NOR4X0 U415 ( .IN1(n295), .IN2(n294), .IN3(n293), .IN4(n292), .QN(N132) );
  XOR2X1 U416 ( .IN1(neighborCount[15]), .IN2(N188), .Q(n304) );
  XOR2X1 U417 ( .IN1(neighborCount[2]), .IN2(N201), .Q(n303) );
  NOR2X0 U418 ( .IN1(n323), .IN2(N203), .QN(n299) );
  OA22X1 U419 ( .IN1(neighborCount[1]), .IN2(n299), .IN3(n299), .IN4(n321), 
        .Q(n302) );
  AND2X1 U420 ( .IN1(N203), .IN2(n323), .Q(n300) );
  OA22X1 U421 ( .IN1(n300), .IN2(n322), .IN3(N202), .IN4(n300), .Q(n301) );
  OR4X1 U422 ( .IN1(n304), .IN2(n303), .IN3(n302), .IN4(n301), .Q(n320) );
  XNOR2X1 U423 ( .IN1(neighborCount[6]), .IN2(N197), .Q(n308) );
  XNOR2X1 U424 ( .IN1(neighborCount[5]), .IN2(N198), .Q(n307) );
  XNOR2X1 U425 ( .IN1(neighborCount[4]), .IN2(N199), .Q(n306) );
  XNOR2X1 U426 ( .IN1(neighborCount[3]), .IN2(N200), .Q(n305) );
  NAND4X0 U427 ( .IN1(n308), .IN2(n307), .IN3(n306), .IN4(n305), .QN(n319) );
  XNOR2X1 U428 ( .IN1(neighborCount[10]), .IN2(N193), .Q(n312) );
  XNOR2X1 U429 ( .IN1(neighborCount[9]), .IN2(N194), .Q(n311) );
  XNOR2X1 U430 ( .IN1(neighborCount[8]), .IN2(N195), .Q(n310) );
  XNOR2X1 U431 ( .IN1(neighborCount[7]), .IN2(N196), .Q(n309) );
  NAND4X0 U432 ( .IN1(n312), .IN2(n311), .IN3(n310), .IN4(n309), .QN(n318) );
  XNOR2X1 U433 ( .IN1(neighborCount[14]), .IN2(N189), .Q(n316) );
  XNOR2X1 U434 ( .IN1(neighborCount[13]), .IN2(N190), .Q(n315) );
  XNOR2X1 U435 ( .IN1(neighborCount[12]), .IN2(N191), .Q(n314) );
  XNOR2X1 U436 ( .IN1(neighborCount[11]), .IN2(N192), .Q(n313) );
  NAND4X0 U437 ( .IN1(n316), .IN2(n315), .IN3(n314), .IN4(n313), .QN(n317) );
  NOR4X0 U438 ( .IN1(n320), .IN2(n319), .IN3(n318), .IN4(n317), .QN(N204) );
endmodule

