`timescale 1ns/1ps
module winnerPolicy_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17;
  wire   [16:0] carry;

  FADDX1 U2_14 ( .A(A[14]), .B(n3), .CI(carry[14]), .CO(carry[15]), .S(
        DIFF[14]) );
  FADDX1 U2_13 ( .A(A[13]), .B(n4), .CI(carry[13]), .CO(carry[14]), .S(
        DIFF[13]) );
  FADDX1 U2_12 ( .A(A[12]), .B(n5), .CI(carry[12]), .CO(carry[13]), .S(
        DIFF[12]) );
  FADDX1 U2_11 ( .A(A[11]), .B(n6), .CI(carry[11]), .CO(carry[12]), .S(
        DIFF[11]) );
  FADDX1 U2_10 ( .A(A[10]), .B(n7), .CI(carry[10]), .CO(carry[11]), .S(
        DIFF[10]) );
  FADDX1 U2_9 ( .A(A[9]), .B(n8), .CI(carry[9]), .CO(carry[10]), .S(DIFF[9])
         );
  FADDX1 U2_8 ( .A(A[8]), .B(n9), .CI(carry[8]), .CO(carry[9]), .S(DIFF[8]) );
  FADDX1 U2_7 ( .A(A[7]), .B(n10), .CI(carry[7]), .CO(carry[8]), .S(DIFF[7])
         );
  FADDX1 U2_6 ( .A(A[6]), .B(n11), .CI(carry[6]), .CO(carry[7]), .S(DIFF[6])
         );
  FADDX1 U2_5 ( .A(A[5]), .B(n12), .CI(carry[5]), .CO(carry[6]), .S(DIFF[5])
         );
  FADDX1 U2_4 ( .A(A[4]), .B(n13), .CI(carry[4]), .CO(carry[5]), .S(DIFF[4])
         );
  FADDX1 U2_3 ( .A(A[3]), .B(n14), .CI(carry[3]), .CO(carry[4]), .S(DIFF[3])
         );
  FADDX1 U2_2 ( .A(A[2]), .B(n15), .CI(carry[2]), .CO(carry[3]), .S(DIFF[2])
         );
  FADDX1 U2_1 ( .A(A[1]), .B(n16), .CI(carry[1]), .CO(carry[2]), .S(DIFF[1])
         );
  XOR3X1 U2_15 ( .IN1(A[15]), .IN2(n2), .IN3(carry[15]), .Q(DIFF[15]) );
  INVX0 U1 ( .INP(B[1]), .ZN(n16) );
  NAND2X1 U2 ( .IN1(B[0]), .IN2(n1), .QN(carry[1]) );
  INVX0 U3 ( .INP(B[2]), .ZN(n15) );
  INVX0 U4 ( .INP(B[3]), .ZN(n14) );
  INVX0 U5 ( .INP(B[4]), .ZN(n13) );
  INVX0 U6 ( .INP(B[5]), .ZN(n12) );
  INVX0 U7 ( .INP(B[6]), .ZN(n11) );
  INVX0 U8 ( .INP(B[7]), .ZN(n10) );
  INVX0 U9 ( .INP(B[8]), .ZN(n9) );
  INVX0 U10 ( .INP(B[9]), .ZN(n8) );
  INVX0 U11 ( .INP(B[10]), .ZN(n7) );
  INVX0 U12 ( .INP(B[11]), .ZN(n6) );
  INVX0 U13 ( .INP(B[12]), .ZN(n5) );
  INVX0 U14 ( .INP(B[13]), .ZN(n4) );
  INVX0 U15 ( .INP(B[14]), .ZN(n3) );
  INVX0 U16 ( .INP(B[15]), .ZN(n2) );
  INVX0 U17 ( .INP(B[0]), .ZN(n17) );
  INVX0 U18 ( .INP(A[0]), .ZN(n1) );
  XOR2X1 U19 ( .IN1(n1), .IN2(n17), .Q(DIFF[0]) );
endmodule


module winnerPolicy_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][5] , \ab[14][5] , \ab[13][5] , \ab[12][5] , \ab[11][5] ,
         \ab[10][5] , \CARRYB[15][5] , \CARRYB[14][5] , \CARRYB[13][5] ,
         \CARRYB[12][5] , \CARRYB[11][5] , n4, n5, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22;
  assign \ab[15][5]  = A[15];
  assign \ab[14][5]  = A[14];
  assign \ab[13][5]  = A[13];
  assign \ab[12][5]  = A[12];
  assign \ab[11][5]  = A[11];
  assign \ab[10][5]  = A[10];

  FADDX1 S4_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(A[5]), .CO(
        \CARRYB[15][5] ), .S(PRODUCT[20]) );
  FADDX1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(A[4]), .CO(
        \CARRYB[14][5] ), .S(PRODUCT[19]) );
  FADDX1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(A[3]), .CO(
        \CARRYB[13][5] ), .S(PRODUCT[18]) );
  FADDX1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(A[2]), .CO(
        \CARRYB[12][5] ), .S(PRODUCT[17]) );
  FADDX1 S2_11_5 ( .A(\ab[11][5] ), .B(n5), .CI(A[1]), .CO(\CARRYB[11][5] ), 
        .S(PRODUCT[16]) );
  AND2X1 U2 ( .IN1(n15), .IN2(\ab[15][5] ), .Q(PRODUCT[31]) );
  OR2X1 U3 ( .IN1(n7), .IN2(A[7]), .Q(n4) );
  NOR2X0 U4 ( .IN1(n14), .IN2(n16), .QN(n15) );
  AND2X1 U5 ( .IN1(\ab[10][5] ), .IN2(A[0]), .Q(n5) );
  AND2X1 U6 ( .IN1(n4), .IN2(n8), .Q(PRODUCT[22]) );
  XNOR2X1 U7 ( .IN1(A[9]), .IN2(n9), .Q(PRODUCT[24]) );
  XNOR2X1 U8 ( .IN1(\ab[10][5] ), .IN2(n10), .Q(PRODUCT[25]) );
  XNOR2X1 U9 ( .IN1(\ab[11][5] ), .IN2(n11), .Q(PRODUCT[26]) );
  XNOR2X1 U10 ( .IN1(\ab[12][5] ), .IN2(n12), .Q(PRODUCT[27]) );
  XNOR2X1 U11 ( .IN1(\ab[13][5] ), .IN2(n13), .Q(PRODUCT[28]) );
  XNOR2X1 U12 ( .IN1(A[8]), .IN2(n8), .Q(PRODUCT[23]) );
  NAND2X1 U13 ( .IN1(n17), .IN2(A[8]), .QN(n9) );
  INVX0 U14 ( .INP(n8), .ZN(n17) );
  NAND2X1 U15 ( .IN1(n22), .IN2(\ab[13][5] ), .QN(n14) );
  INVX0 U16 ( .INP(n13), .ZN(n22) );
  NAND2X1 U17 ( .IN1(n19), .IN2(\ab[10][5] ), .QN(n11) );
  INVX0 U18 ( .INP(n10), .ZN(n19) );
  NAND2X1 U19 ( .IN1(n21), .IN2(\ab[12][5] ), .QN(n13) );
  INVX0 U20 ( .INP(n12), .ZN(n21) );
  NAND2X1 U21 ( .IN1(n18), .IN2(A[9]), .QN(n10) );
  INVX0 U22 ( .INP(n9), .ZN(n18) );
  NAND2X1 U23 ( .IN1(n20), .IN2(\ab[11][5] ), .QN(n12) );
  INVX0 U24 ( .INP(n11), .ZN(n20) );
  AND2X1 U25 ( .IN1(A[6]), .IN2(\CARRYB[15][5] ), .Q(n7) );
  INVX0 U26 ( .INP(\ab[14][5] ), .ZN(n16) );
  XOR2X1 U27 ( .IN1(\CARRYB[15][5] ), .IN2(A[6]), .Q(PRODUCT[21]) );
  XOR2X1 U28 ( .IN1(A[0]), .IN2(\ab[10][5] ), .Q(PRODUCT[15]) );
  NAND2X0 U29 ( .IN1(n7), .IN2(A[7]), .QN(n8) );
  XOR2X1 U30 ( .IN1(n16), .IN2(n14), .Q(PRODUCT[29]) );
  XOR2X1 U31 ( .IN1(\ab[15][5] ), .IN2(n15), .Q(PRODUCT[30]) );
endmodule


module winnerPolicy_DW01_add_2 ( A, B, CI, SUM, CO );
  input [29:0] A;
  input [29:0] B;
  output [29:0] SUM;
  input CI;
  output CO;
  wire   \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] , \A[7] ,
         \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1, n2, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n56, n57;
  assign SUM[15] = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  OR2X1 U2 ( .IN1(B[16]), .IN2(A[16]), .Q(n1) );
  NAND2X1 U3 ( .IN1(n10), .IN2(A[21]), .QN(n37) );
  INVX0 U4 ( .INP(n41), .ZN(n10) );
  XOR2X1 U5 ( .IN1(B[29]), .IN2(n2), .Q(SUM[29]) );
  AO22X1 U6 ( .IN1(n15), .IN2(B[28]), .IN3(n16), .IN4(A[28]), .Q(n2) );
  INVX0 U7 ( .INP(n18), .ZN(n4) );
  INVX0 U8 ( .INP(n43), .ZN(n11) );
  INVX0 U9 ( .INP(n22), .ZN(n5) );
  INVX0 U10 ( .INP(n26), .ZN(n6) );
  INVX0 U11 ( .INP(n30), .ZN(n7) );
  INVX0 U12 ( .INP(n34), .ZN(n8) );
  INVX0 U13 ( .INP(n38), .ZN(n9) );
  INVX0 U14 ( .INP(n47), .ZN(n12) );
  INVX0 U15 ( .INP(n51), .ZN(n13) );
  XNOR2X1 U16 ( .IN1(A[21]), .IN2(n41), .Q(SUM[21]) );
  AND2X1 U17 ( .IN1(n1), .IN2(n54), .Q(SUM[16]) );
  INVX0 U18 ( .INP(n55), .ZN(n14) );
  OR2X1 U19 ( .IN1(A[28]), .IN2(n16), .Q(n15) );
  XOR3X1 U20 ( .IN1(B[28]), .IN2(A[28]), .IN3(n16), .Q(SUM[28]) );
  OAI21X1 U21 ( .IN1(n17), .IN2(n18), .IN3(n19), .QN(n16) );
  XOR2X1 U22 ( .IN1(n20), .IN2(n17), .Q(SUM[27]) );
  OA21X1 U23 ( .IN1(n21), .IN2(n22), .IN3(n23), .Q(n17) );
  NAND2X0 U24 ( .IN1(n4), .IN2(n19), .QN(n20) );
  NAND2X0 U25 ( .IN1(B[27]), .IN2(A[27]), .QN(n19) );
  NOR2X0 U26 ( .IN1(B[27]), .IN2(A[27]), .QN(n18) );
  XOR2X1 U27 ( .IN1(n24), .IN2(n21), .Q(SUM[26]) );
  OA21X1 U28 ( .IN1(n25), .IN2(n26), .IN3(n27), .Q(n21) );
  NAND2X0 U29 ( .IN1(n5), .IN2(n23), .QN(n24) );
  NAND2X0 U30 ( .IN1(B[26]), .IN2(A[26]), .QN(n23) );
  NOR2X0 U31 ( .IN1(B[26]), .IN2(A[26]), .QN(n22) );
  XOR2X1 U32 ( .IN1(n28), .IN2(n25), .Q(SUM[25]) );
  OA21X1 U33 ( .IN1(n29), .IN2(n30), .IN3(n31), .Q(n25) );
  NAND2X0 U34 ( .IN1(n6), .IN2(n27), .QN(n28) );
  NAND2X0 U35 ( .IN1(B[25]), .IN2(A[25]), .QN(n27) );
  NOR2X0 U36 ( .IN1(B[25]), .IN2(A[25]), .QN(n26) );
  XOR2X1 U37 ( .IN1(n32), .IN2(n29), .Q(SUM[24]) );
  OA21X1 U38 ( .IN1(n33), .IN2(n34), .IN3(n35), .Q(n29) );
  NAND2X0 U39 ( .IN1(n7), .IN2(n31), .QN(n32) );
  NAND2X0 U40 ( .IN1(B[24]), .IN2(A[24]), .QN(n31) );
  NOR2X0 U41 ( .IN1(B[24]), .IN2(A[24]), .QN(n30) );
  XOR2X1 U42 ( .IN1(n36), .IN2(n33), .Q(SUM[23]) );
  OA21X1 U43 ( .IN1(n37), .IN2(n38), .IN3(n39), .Q(n33) );
  NAND2X0 U44 ( .IN1(n8), .IN2(n35), .QN(n36) );
  NAND2X0 U45 ( .IN1(B[23]), .IN2(A[23]), .QN(n35) );
  NOR2X0 U46 ( .IN1(B[23]), .IN2(A[23]), .QN(n34) );
  XOR2X1 U47 ( .IN1(n40), .IN2(n37), .Q(SUM[22]) );
  NAND2X0 U48 ( .IN1(n9), .IN2(n39), .QN(n40) );
  NAND2X0 U49 ( .IN1(B[22]), .IN2(A[22]), .QN(n39) );
  NOR2X0 U50 ( .IN1(B[22]), .IN2(A[22]), .QN(n38) );
  OA21X1 U51 ( .IN1(n42), .IN2(n43), .IN3(n44), .Q(n41) );
  XOR2X1 U52 ( .IN1(n45), .IN2(n42), .Q(SUM[20]) );
  OA21X1 U53 ( .IN1(n46), .IN2(n47), .IN3(n48), .Q(n42) );
  NAND2X0 U54 ( .IN1(n11), .IN2(n44), .QN(n45) );
  NAND2X0 U55 ( .IN1(B[20]), .IN2(A[20]), .QN(n44) );
  NOR2X0 U56 ( .IN1(B[20]), .IN2(A[20]), .QN(n43) );
  XOR2X1 U57 ( .IN1(n49), .IN2(n46), .Q(SUM[19]) );
  OA21X1 U58 ( .IN1(n50), .IN2(n51), .IN3(n52), .Q(n46) );
  NAND2X0 U59 ( .IN1(n12), .IN2(n48), .QN(n49) );
  NAND2X0 U60 ( .IN1(B[19]), .IN2(A[19]), .QN(n48) );
  NOR2X0 U61 ( .IN1(B[19]), .IN2(A[19]), .QN(n47) );
  XOR2X1 U62 ( .IN1(n53), .IN2(n50), .Q(SUM[18]) );
  OA21X1 U63 ( .IN1(n54), .IN2(n55), .IN3(n56), .Q(n50) );
  NAND2X0 U64 ( .IN1(n13), .IN2(n52), .QN(n53) );
  NAND2X0 U65 ( .IN1(B[18]), .IN2(A[18]), .QN(n52) );
  NOR2X0 U66 ( .IN1(B[18]), .IN2(A[18]), .QN(n51) );
  XOR2X1 U67 ( .IN1(n57), .IN2(n54), .Q(SUM[17]) );
  NAND2X0 U68 ( .IN1(n14), .IN2(n56), .QN(n57) );
  NAND2X0 U69 ( .IN1(B[17]), .IN2(A[17]), .QN(n56) );
  NOR2X0 U70 ( .IN1(B[17]), .IN2(A[17]), .QN(n55) );
  NAND2X0 U71 ( .IN1(B[16]), .IN2(A[16]), .QN(n54) );
endmodule


module winnerPolicy_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [15:0] A;
  input [15:0] B;
  output [31:0] PRODUCT;
  input TC;
  wire   \ab[15][9] , \ab[14][9] , \ab[13][9] , \ab[12][9] , \ab[11][9] ,
         \ab[10][9] , \ab[9][9] , \ab[8][9] , \ab[7][9] , \ab[6][9] ,
         \ab[5][9] , \ab[4][9] , \ab[3][9] , \ab[2][9] , \ab[1][9] ,
         \ab[0][9] , \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][5] , \CARRYB[15][4] , \CARRYB[15][3] ,
         \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][5] , \CARRYB[14][4] ,
         \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] , \CARRYB[13][14] ,
         \CARRYB[13][13] , \CARRYB[13][12] , \CARRYB[13][11] ,
         \CARRYB[13][10] , \CARRYB[13][9] , \CARRYB[13][8] , \CARRYB[13][7] ,
         \CARRYB[13][5] , \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] ,
         \CARRYB[13][1] , \CARRYB[12][14] , \CARRYB[12][13] , \CARRYB[12][12] ,
         \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] , \CARRYB[12][8] ,
         \CARRYB[12][7] , \CARRYB[12][5] , \CARRYB[12][4] , \CARRYB[12][3] ,
         \CARRYB[12][2] , \CARRYB[12][1] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][5] , \CARRYB[11][4] ,
         \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] , \CARRYB[10][14] ,
         \CARRYB[10][13] , \CARRYB[10][12] , \CARRYB[10][11] ,
         \CARRYB[10][10] , \CARRYB[10][9] , \CARRYB[10][8] , \CARRYB[10][7] ,
         \CARRYB[10][5] , \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] ,
         \CARRYB[10][1] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][5] , \CARRYB[9][4] , \CARRYB[9][3] ,
         \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][5] , \CARRYB[8][4] ,
         \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[6][14] , \CARRYB[6][13] , \CARRYB[6][12] , \CARRYB[6][11] ,
         \CARRYB[6][10] , \CARRYB[6][9] , \CARRYB[6][8] , \CARRYB[6][7] ,
         \CARRYB[6][5] , \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] ,
         \CARRYB[6][1] , \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] ,
         \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] ,
         \CARRYB[5][7] , \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] ,
         \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[4][14] , \CARRYB[4][13] ,
         \CARRYB[4][12] , \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] ,
         \CARRYB[4][8] , \CARRYB[4][7] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][5] ,
         \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] , \CARRYB[3][1] ,
         \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] , \CARRYB[2][11] ,
         \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] , \CARRYB[2][7] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][3] ,
         \CARRYB[1][2] , \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] ,
         \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] ,
         \SUMB[15][7] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][5] , \SUMB[14][4] ,
         \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][14] ,
         \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] ,
         \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] ,
         \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] ,
         \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] ,
         \SUMB[12][1] , \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] ,
         \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] ,
         \SUMB[11][7] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][5] , \SUMB[10][4] ,
         \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][14] ,
         \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] ,
         \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][5] , \SUMB[8][4] ,
         \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][5] , \SUMB[7][4] ,
         \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][14] ,
         \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] , \SUMB[6][10] ,
         \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][5] , \SUMB[6][4] ,
         \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] , \SUMB[5][14] ,
         \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] , \SUMB[5][10] ,
         \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][5] , \SUMB[5][4] ,
         \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][14] ,
         \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] , \SUMB[4][10] ,
         \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][5] , \SUMB[4][4] ,
         \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][5] , \SUMB[3][4] ,
         \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][14] ,
         \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] ,
         \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][4] , \SUMB[1][3] ,
         \SUMB[1][2] , \SUMB[1][1] , \A1[28] , \A1[27] , \A1[26] , \A1[25] ,
         \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[19] , \A1[18] , \A1[17] ,
         \A1[16] , \A1[15] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23;
  assign \ab[15][9]  = A[15];
  assign \ab[14][9]  = A[14];
  assign \ab[13][9]  = A[13];
  assign \ab[12][9]  = A[12];
  assign \ab[11][9]  = A[11];
  assign \ab[10][9]  = A[10];
  assign \ab[9][9]  = A[9];
  assign \ab[8][9]  = A[8];
  assign \ab[7][9]  = A[7];
  assign \ab[6][9]  = A[6];
  assign \ab[5][9]  = A[5];
  assign \ab[4][9]  = A[4];
  assign \ab[3][9]  = A[3];
  assign \ab[2][9]  = A[2];
  assign \ab[1][9]  = A[1];
  assign PRODUCT[1] = \ab[0][9] ;
  assign \ab[0][9]  = A[0];

  FADDX1 S4_1 ( .A(\ab[15][9] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), .CO(
        \CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FADDX1 S4_2 ( .A(\ab[15][9] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), .CO(
        \CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FADDX1 S4_3 ( .A(\ab[15][9] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), .CO(
        \CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FADDX1 S4_4 ( .A(\ab[15][9] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), .CO(
        \CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FADDX1 S4_5 ( .A(\ab[15][9] ), .B(\CARRYB[14][5] ), .CI(\SUMB[13][7] ), .CO(
        \CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FADDX1 S4_7 ( .A(\ab[15][9] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), .CO(
        \CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FADDX1 S4_8 ( .A(\ab[15][9] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), .CO(
        \CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FADDX1 S4_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FADDX1 S4_10 ( .A(\ab[15][9] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FADDX1 S4_11 ( .A(\ab[15][9] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FADDX1 S4_12 ( .A(\ab[15][9] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FADDX1 S4_13 ( .A(\ab[15][9] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FADDX1 S5_14 ( .A(\ab[15][9] ), .B(\CARRYB[14][14] ), .CI(\ab[14][9] ), .CO(
        \CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FADDX1 S2_14_1 ( .A(\ab[14][9] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FADDX1 S2_14_2 ( .A(\ab[14][9] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FADDX1 S2_14_3 ( .A(\ab[14][9] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FADDX1 S2_14_4 ( .A(\ab[14][9] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FADDX1 S2_14_5 ( .A(\ab[14][9] ), .B(\CARRYB[13][5] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FADDX1 S2_14_7 ( .A(\ab[14][9] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FADDX1 S2_14_8 ( .A(\ab[14][9] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FADDX1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FADDX1 S2_14_10 ( .A(\ab[14][9] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FADDX1 S2_14_11 ( .A(\ab[14][9] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FADDX1 S2_14_12 ( .A(\ab[14][9] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FADDX1 S2_14_13 ( .A(\ab[14][9] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FADDX1 S3_14_14 ( .A(\ab[14][9] ), .B(\CARRYB[13][14] ), .CI(\ab[13][9] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FADDX1 S2_13_1 ( .A(\ab[13][9] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FADDX1 S2_13_2 ( .A(\ab[13][9] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FADDX1 S2_13_3 ( .A(\ab[13][9] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FADDX1 S2_13_4 ( .A(\ab[13][9] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FADDX1 S2_13_5 ( .A(\ab[13][9] ), .B(\CARRYB[12][5] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FADDX1 S2_13_7 ( .A(\ab[13][9] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FADDX1 S2_13_8 ( .A(\ab[13][9] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FADDX1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FADDX1 S2_13_10 ( .A(\ab[13][9] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FADDX1 S2_13_11 ( .A(\ab[13][9] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FADDX1 S2_13_12 ( .A(\ab[13][9] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FADDX1 S2_13_13 ( .A(\ab[13][9] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FADDX1 S3_13_14 ( .A(\ab[13][9] ), .B(\CARRYB[12][14] ), .CI(\ab[12][9] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FADDX1 S2_12_1 ( .A(\ab[12][9] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FADDX1 S2_12_2 ( .A(\ab[12][9] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FADDX1 S2_12_3 ( .A(\ab[12][9] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FADDX1 S2_12_4 ( .A(\ab[12][9] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FADDX1 S2_12_5 ( .A(\ab[12][9] ), .B(\CARRYB[11][5] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FADDX1 S2_12_7 ( .A(\ab[12][9] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FADDX1 S2_12_8 ( .A(\ab[12][9] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FADDX1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FADDX1 S2_12_10 ( .A(\ab[12][9] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FADDX1 S2_12_11 ( .A(\ab[12][9] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FADDX1 S2_12_12 ( .A(\ab[12][9] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FADDX1 S2_12_13 ( .A(\ab[12][9] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FADDX1 S3_12_14 ( .A(\ab[12][9] ), .B(\CARRYB[11][14] ), .CI(\ab[11][9] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FADDX1 S2_11_1 ( .A(\ab[11][9] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FADDX1 S2_11_2 ( .A(\ab[11][9] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FADDX1 S2_11_3 ( .A(\ab[11][9] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FADDX1 S2_11_4 ( .A(\ab[11][9] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FADDX1 S2_11_5 ( .A(\ab[11][9] ), .B(\CARRYB[10][5] ), .CI(\SUMB[9][7] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FADDX1 S2_11_7 ( .A(\ab[11][9] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FADDX1 S2_11_8 ( .A(\ab[11][9] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FADDX1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FADDX1 S2_11_10 ( .A(\ab[11][9] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FADDX1 S2_11_11 ( .A(\ab[11][9] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FADDX1 S2_11_12 ( .A(\ab[11][9] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FADDX1 S2_11_13 ( .A(\ab[11][9] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FADDX1 S3_11_14 ( .A(\ab[11][9] ), .B(\CARRYB[10][14] ), .CI(\ab[10][9] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FADDX1 S2_10_1 ( .A(\ab[10][9] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), 
        .CO(\CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FADDX1 S2_10_2 ( .A(\ab[10][9] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), 
        .CO(\CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FADDX1 S2_10_3 ( .A(\ab[10][9] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), 
        .CO(\CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FADDX1 S2_10_4 ( .A(\ab[10][9] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), 
        .CO(\CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FADDX1 S2_10_5 ( .A(\ab[10][9] ), .B(\CARRYB[9][5] ), .CI(\SUMB[8][7] ), 
        .CO(\CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FADDX1 S2_10_7 ( .A(\ab[10][9] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), 
        .CO(\CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FADDX1 S2_10_8 ( .A(\ab[10][9] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), 
        .CO(\CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FADDX1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FADDX1 S2_10_10 ( .A(\ab[10][9] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FADDX1 S2_10_11 ( .A(\ab[10][9] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FADDX1 S2_10_12 ( .A(\ab[10][9] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FADDX1 S2_10_13 ( .A(\ab[10][9] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FADDX1 S3_10_14 ( .A(\ab[10][9] ), .B(\CARRYB[9][14] ), .CI(\ab[9][9] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FADDX1 S2_9_1 ( .A(\ab[9][9] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FADDX1 S2_9_2 ( .A(\ab[9][9] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FADDX1 S2_9_3 ( .A(\ab[9][9] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FADDX1 S2_9_4 ( .A(\ab[9][9] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FADDX1 S2_9_5 ( .A(\ab[9][9] ), .B(\CARRYB[8][5] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FADDX1 S2_9_7 ( .A(\ab[9][9] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FADDX1 S2_9_8 ( .A(\ab[9][9] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FADDX1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FADDX1 S2_9_10 ( .A(\ab[9][9] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FADDX1 S2_9_11 ( .A(\ab[9][9] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FADDX1 S2_9_12 ( .A(\ab[9][9] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FADDX1 S2_9_13 ( .A(\ab[9][9] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FADDX1 S3_9_14 ( .A(\ab[9][9] ), .B(\CARRYB[8][14] ), .CI(\ab[8][9] ), .CO(
        \CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FADDX1 S2_8_1 ( .A(\ab[8][9] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FADDX1 S2_8_2 ( .A(\ab[8][9] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FADDX1 S2_8_3 ( .A(\ab[8][9] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FADDX1 S2_8_4 ( .A(\ab[8][9] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FADDX1 S2_8_5 ( .A(\ab[8][9] ), .B(\CARRYB[7][5] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FADDX1 S2_8_7 ( .A(\ab[8][9] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FADDX1 S2_8_8 ( .A(\ab[8][9] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FADDX1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FADDX1 S2_8_10 ( .A(\ab[8][9] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FADDX1 S2_8_11 ( .A(\ab[8][9] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FADDX1 S2_8_12 ( .A(\ab[8][9] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FADDX1 S2_8_13 ( .A(\ab[8][9] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FADDX1 S3_8_14 ( .A(\ab[8][9] ), .B(\CARRYB[7][14] ), .CI(\ab[7][9] ), .CO(
        \CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FADDX1 S2_7_1 ( .A(\ab[7][9] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FADDX1 S2_7_2 ( .A(\ab[7][9] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FADDX1 S2_7_3 ( .A(\ab[7][9] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FADDX1 S2_7_4 ( .A(\ab[7][9] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FADDX1 S2_7_5 ( .A(\ab[7][9] ), .B(\CARRYB[6][5] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FADDX1 S2_7_7 ( .A(\ab[7][9] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FADDX1 S2_7_8 ( .A(\ab[7][9] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FADDX1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FADDX1 S2_7_10 ( .A(\ab[7][9] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FADDX1 S2_7_11 ( .A(\ab[7][9] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FADDX1 S2_7_12 ( .A(\ab[7][9] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FADDX1 S2_7_13 ( .A(\ab[7][9] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FADDX1 S3_7_14 ( .A(\ab[7][9] ), .B(\CARRYB[6][14] ), .CI(\ab[6][9] ), .CO(
        \CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FADDX1 S2_6_1 ( .A(\ab[6][9] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FADDX1 S2_6_2 ( .A(\ab[6][9] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FADDX1 S2_6_3 ( .A(\ab[6][9] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FADDX1 S2_6_4 ( .A(\ab[6][9] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FADDX1 S2_6_5 ( .A(\ab[6][9] ), .B(\CARRYB[5][5] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FADDX1 S2_6_7 ( .A(\ab[6][9] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FADDX1 S2_6_8 ( .A(\ab[6][9] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FADDX1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FADDX1 S2_6_10 ( .A(\ab[6][9] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FADDX1 S2_6_11 ( .A(\ab[6][9] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FADDX1 S2_6_12 ( .A(\ab[6][9] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FADDX1 S2_6_13 ( .A(\ab[6][9] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FADDX1 S3_6_14 ( .A(\ab[6][9] ), .B(\CARRYB[5][14] ), .CI(\ab[5][9] ), .CO(
        \CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FADDX1 S2_5_1 ( .A(\ab[5][9] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FADDX1 S2_5_2 ( .A(\ab[5][9] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FADDX1 S2_5_3 ( .A(\ab[5][9] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FADDX1 S2_5_4 ( .A(\ab[5][9] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FADDX1 S2_5_5 ( .A(\ab[5][9] ), .B(\CARRYB[4][5] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FADDX1 S2_5_7 ( .A(\ab[5][9] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FADDX1 S2_5_8 ( .A(\ab[5][9] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FADDX1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FADDX1 S2_5_10 ( .A(\ab[5][9] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FADDX1 S2_5_11 ( .A(\ab[5][9] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FADDX1 S2_5_12 ( .A(\ab[5][9] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FADDX1 S2_5_13 ( .A(\ab[5][9] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FADDX1 S3_5_14 ( .A(\ab[5][9] ), .B(\CARRYB[4][14] ), .CI(\ab[4][9] ), .CO(
        \CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FADDX1 S2_4_1 ( .A(\ab[4][9] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FADDX1 S2_4_2 ( .A(\ab[4][9] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FADDX1 S2_4_3 ( .A(\ab[4][9] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FADDX1 S2_4_4 ( .A(\ab[4][9] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FADDX1 S2_4_5 ( .A(\ab[4][9] ), .B(\CARRYB[3][5] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FADDX1 S2_4_7 ( .A(\ab[4][9] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FADDX1 S2_4_8 ( .A(\ab[4][9] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FADDX1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FADDX1 S2_4_10 ( .A(\ab[4][9] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FADDX1 S2_4_11 ( .A(\ab[4][9] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FADDX1 S2_4_12 ( .A(\ab[4][9] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FADDX1 S2_4_13 ( .A(\ab[4][9] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FADDX1 S3_4_14 ( .A(\ab[4][9] ), .B(\CARRYB[3][14] ), .CI(\ab[3][9] ), .CO(
        \CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FADDX1 S2_3_1 ( .A(\ab[3][9] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FADDX1 S2_3_2 ( .A(\ab[3][9] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FADDX1 S2_3_3 ( .A(\ab[3][9] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FADDX1 S2_3_4 ( .A(\ab[3][9] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FADDX1 S2_3_5 ( .A(\ab[3][9] ), .B(n3), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FADDX1 S2_3_7 ( .A(\ab[3][9] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FADDX1 S2_3_8 ( .A(\ab[3][9] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FADDX1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FADDX1 S2_3_10 ( .A(\ab[3][9] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FADDX1 S2_3_11 ( .A(\ab[3][9] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FADDX1 S2_3_12 ( .A(\ab[3][9] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FADDX1 S2_3_13 ( .A(\ab[3][9] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FADDX1 S3_3_14 ( .A(\ab[3][9] ), .B(\CARRYB[2][14] ), .CI(\ab[2][9] ), .CO(
        \CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FADDX1 S2_2_1 ( .A(\ab[2][9] ), .B(n17), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FADDX1 S2_2_2 ( .A(\ab[2][9] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FADDX1 S2_2_3 ( .A(\ab[2][9] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FADDX1 S2_2_4 ( .A(\ab[2][9] ), .B(n16), .CI(\ab[1][9] ), .CO(\CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FADDX1 S2_2_7 ( .A(\ab[2][9] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FADDX1 S2_2_8 ( .A(\ab[2][9] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FADDX1 S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][10] ), 
        .CO(\CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FADDX1 S2_2_10 ( .A(\ab[2][9] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FADDX1 S2_2_11 ( .A(\ab[2][9] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FADDX1 S2_2_12 ( .A(\ab[2][9] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FADDX1 S2_2_13 ( .A(\ab[2][9] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FADDX1 S3_2_14 ( .A(\ab[2][9] ), .B(n17), .CI(\ab[1][9] ), .CO(
        \CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  winnerPolicy_DW01_add_2 FS_1 ( .A({1'b0, \A1[28] , \A1[27] , \A1[26] , 
        \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \SUMB[15][7] , 
        \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \SUMB[15][1] , 
        \SUMB[14][1] , \SUMB[13][1] , \SUMB[12][1] , \SUMB[11][1] , 
        \SUMB[10][1] , \SUMB[9][1] , \SUMB[8][1] , \SUMB[7][1] , \SUMB[6][1] , 
        \SUMB[5][1] , \SUMB[4][1] , \SUMB[3][1] , \SUMB[2][1] , \SUMB[1][1] }), 
        .B({n18, n15, n6, n7, n8, n9, n10, n11, 1'b0, n12, n13, n14, n4, n5, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[31:2]) );
  AND2X1 U2 ( .IN1(\ab[2][9] ), .IN2(\ab[0][9] ), .Q(n3) );
  AND2X1 U3 ( .IN1(\CARRYB[15][2] ), .IN2(\SUMB[15][3] ), .Q(n4) );
  AND2X1 U4 ( .IN1(\CARRYB[15][1] ), .IN2(\SUMB[15][2] ), .Q(n5) );
  AND2X1 U5 ( .IN1(\CARRYB[15][12] ), .IN2(\SUMB[15][13] ), .Q(n6) );
  AND2X1 U6 ( .IN1(\CARRYB[15][11] ), .IN2(\SUMB[15][12] ), .Q(n7) );
  AND2X1 U7 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .Q(n8) );
  AND2X1 U8 ( .IN1(\CARRYB[15][9] ), .IN2(\SUMB[15][10] ), .Q(n9) );
  AND2X1 U9 ( .IN1(\CARRYB[15][8] ), .IN2(\SUMB[15][9] ), .Q(n10) );
  AND2X1 U10 ( .IN1(\CARRYB[15][7] ), .IN2(\SUMB[15][8] ), .Q(n11) );
  AND2X1 U11 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[14][7] ), .Q(n12) );
  AND2X1 U12 ( .IN1(\CARRYB[15][4] ), .IN2(\SUMB[15][5] ), .Q(n13) );
  AND2X1 U13 ( .IN1(\CARRYB[15][3] ), .IN2(\SUMB[15][4] ), .Q(n14) );
  AND2X1 U14 ( .IN1(\CARRYB[15][13] ), .IN2(\SUMB[15][14] ), .Q(n15) );
  INVX0 U15 ( .INP(n19), .ZN(\CARRYB[1][2] ) );
  NAND2X1 U16 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .QN(n19) );
  INVX0 U17 ( .INP(n20), .ZN(\CARRYB[1][3] ) );
  NAND2X1 U18 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .QN(n20) );
  AND2X1 U19 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .Q(n16) );
  INVX0 U20 ( .INP(n21), .ZN(\CARRYB[1][11] ) );
  NAND2X1 U21 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .QN(n21) );
  INVX0 U22 ( .INP(n22), .ZN(\CARRYB[1][12] ) );
  NAND2X1 U23 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .QN(n22) );
  INVX0 U24 ( .INP(n23), .ZN(\CARRYB[1][13] ) );
  NAND2X1 U25 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .QN(n23) );
  AND2X1 U26 ( .IN1(\ab[0][9] ), .IN2(\ab[1][9] ), .Q(n17) );
  AND2X1 U27 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[15][9] ), .Q(n18) );
  XOR2X1 U28 ( .IN1(\CARRYB[15][1] ), .IN2(\SUMB[15][2] ), .Q(\A1[15] ) );
  XOR2X1 U29 ( .IN1(\CARRYB[15][2] ), .IN2(\SUMB[15][3] ), .Q(\A1[16] ) );
  XOR2X1 U30 ( .IN1(\CARRYB[15][3] ), .IN2(\SUMB[15][4] ), .Q(\A1[17] ) );
  XOR2X1 U31 ( .IN1(\CARRYB[15][4] ), .IN2(\SUMB[15][5] ), .Q(\A1[18] ) );
  XOR2X1 U32 ( .IN1(\CARRYB[15][5] ), .IN2(\SUMB[14][7] ), .Q(\A1[19] ) );
  XOR2X1 U33 ( .IN1(\CARRYB[15][7] ), .IN2(\SUMB[15][8] ), .Q(\A1[21] ) );
  XOR2X1 U34 ( .IN1(\CARRYB[15][8] ), .IN2(\SUMB[15][9] ), .Q(\A1[22] ) );
  XOR2X1 U35 ( .IN1(\CARRYB[15][9] ), .IN2(\SUMB[15][10] ), .Q(\A1[23] ) );
  XOR2X1 U36 ( .IN1(\CARRYB[15][10] ), .IN2(\SUMB[15][11] ), .Q(\A1[24] ) );
  XOR2X1 U37 ( .IN1(\CARRYB[15][11] ), .IN2(\SUMB[15][12] ), .Q(\A1[25] ) );
  XOR2X1 U38 ( .IN1(\CARRYB[15][12] ), .IN2(\SUMB[15][13] ), .Q(\A1[26] ) );
  XOR2X1 U39 ( .IN1(\CARRYB[15][13] ), .IN2(\SUMB[15][14] ), .Q(\A1[27] ) );
  XOR2X1 U40 ( .IN1(\CARRYB[15][14] ), .IN2(\ab[15][9] ), .Q(\A1[28] ) );
  XOR2X1 U41 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][1] ) );
  XOR2X1 U42 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][2] ) );
  XOR2X1 U43 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][3] ) );
  XOR2X1 U44 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][4] ) );
  XOR2X1 U45 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][7] ) );
  XOR2X1 U46 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][8] ) );
  XOR2X1 U47 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][9] ) );
  XOR2X1 U48 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][10] ) );
  XOR2X1 U49 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][11] ) );
  XOR2X1 U50 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][12] ) );
  XOR2X1 U51 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][13] ) );
  XOR2X1 U52 ( .IN1(\ab[1][9] ), .IN2(\ab[0][9] ), .Q(\SUMB[1][14] ) );
  XOR2X1 U53 ( .IN1(\ab[0][9] ), .IN2(\ab[2][9] ), .Q(\SUMB[2][5] ) );
endmodule


module winnerPolicy ( clock, nrst, en, start_winnerPolicy, mybest, besthop, 
        bestvalue, bestneighborID, MY_NODE_ID, address, data_in, wr_en, 
        data_out, epsilon_step, nexthop, done_winnerPolicy, en_rng, rng_out, 
        rng_out_4bit, rng_address, start_rngAddress, done_rng_address, 
        betterNeighborCount, which );
  input [15:0] mybest;
  input [15:0] besthop;
  input [15:0] bestvalue;
  input [15:0] bestneighborID;
  input [15:0] MY_NODE_ID;
  output [10:0] address;
  input [15:0] data_in;
  output [15:0] data_out;
  input [15:0] epsilon_step;
  output [15:0] nexthop;
  input [15:0] rng_out;
  input [15:0] rng_out_4bit;
  input [15:0] rng_address;
  output [15:0] betterNeighborCount;
  output [15:0] which;
  input clock, nrst, en, start_winnerPolicy, done_rng_address;
  output wr_en, done_winnerPolicy, en_rng, start_rngAddress;
  wire   one, two, three, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N165, N166, N167, N168, N169,
         N170, N171, N172, N173, N174, N175, N176, N177, N178, N179, N180,
         N181, N182, N183, N184, N185, N186, N187, N188, N189, N190, N191,
         N192, N193, N194, N195, N196, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N476, N477, N478, N479, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, N229, N228, N227,
         N226, N225, N224, N223, N222, N221, N220, N219, N218, N217, N216,
         N215, N214, N213, \add_121/carry[10] , \add_121/carry[9] ,
         \add_121/carry[8] , \add_121/carry[7] , \add_121/carry[6] ,
         \add_121/carry[5] , \add_173/carry[31] , \add_173/carry[30] ,
         \add_173/carry[29] , \add_173/carry[28] , \add_173/carry[27] ,
         \add_173/carry[26] , \add_173/carry[25] , \add_173/carry[24] ,
         \add_173/carry[23] , \add_173/carry[22] , \add_173/carry[21] ,
         \add_173/carry[20] , \add_173/carry[19] , \add_173/carry[18] ,
         \add_173/carry[17] , \add_173/carry[16] , n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595;
  wire   [3:0] state;
  wire   [15:0] epsilon_buf;
  wire   [31:0] _left;
  wire   [31:0] _right3;
  wire   [31:0] _right;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;
  assign N119 = rng_address[0];
  assign N120 = rng_address[1];
  assign N235 = mybest[0];
  assign N236 = mybest[1];
  assign N237 = mybest[2];
  assign N238 = mybest[3];
  assign N239 = mybest[4];
  assign N240 = mybest[5];
  assign N241 = mybest[6];
  assign N242 = mybest[7];
  assign N243 = mybest[8];
  assign N244 = mybest[9];

  DFFX1 \_right_reg[7]  ( .D(n201), .CLK(clock), .Q(_right[7]) );
  DFFX1 \_right_reg[8]  ( .D(n200), .CLK(clock), .Q(_right[8]) );
  DFFX1 \_right_reg[9]  ( .D(n199), .CLK(clock), .Q(_right[9]) );
  DFFX1 \_right_reg[10]  ( .D(n198), .CLK(clock), .Q(_right[10]) );
  DFFX1 \_right_reg[11]  ( .D(n197), .CLK(clock), .Q(_right[11]) );
  DFFX1 \_right_reg[12]  ( .D(n196), .CLK(clock), .Q(_right[12]) );
  DFFX1 \_right_reg[13]  ( .D(n195), .CLK(clock), .Q(_right[13]) );
  DFFX1 \_right_reg[14]  ( .D(n194), .CLK(clock), .Q(_right[14]) );
  DFFX1 \_right_reg[15]  ( .D(n193), .CLK(clock), .Q(_right[15]) );
  DFFX1 \_right_reg[16]  ( .D(n192), .CLK(clock), .Q(_right[16]) );
  DFFX1 \_right_reg[17]  ( .D(n191), .CLK(clock), .Q(_right[17]) );
  DFFX1 \_right_reg[18]  ( .D(n190), .CLK(clock), .Q(_right[18]) );
  DFFX1 \_right_reg[19]  ( .D(n189), .CLK(clock), .Q(_right[19]) );
  DFFX1 \_right_reg[20]  ( .D(n188), .CLK(clock), .Q(_right[20]) );
  DFFX1 \_right_reg[21]  ( .D(n187), .CLK(clock), .Q(_right[21]) );
  DFFX1 \_right_reg[22]  ( .D(n186), .CLK(clock), .Q(_right[22]) );
  DFFX1 \_right_reg[23]  ( .D(n185), .CLK(clock), .Q(_right[23]) );
  DFFX1 \_right_reg[24]  ( .D(n184), .CLK(clock), .Q(_right[24]) );
  DFFX1 \_right_reg[25]  ( .D(n183), .CLK(clock), .Q(_right[25]) );
  DFFX1 \_right_reg[26]  ( .D(n182), .CLK(clock), .Q(_right[26]) );
  DFFX1 \_right_reg[27]  ( .D(n181), .CLK(clock), .Q(_right[27]) );
  DFFX1 \_right_reg[28]  ( .D(n180), .CLK(clock), .Q(_right[28]) );
  DFFX1 \_right_reg[29]  ( .D(n179), .CLK(clock), .Q(_right[29]) );
  DFFX1 \_right_reg[30]  ( .D(n178), .CLK(clock), .Q(_right[30]) );
  DFFX1 \_right_reg[31]  ( .D(n177), .CLK(clock), .Q(_right[31]) );
  DFFX1 \_right3_reg[31]  ( .D(n144), .CLK(clock), .Q(_right3[31]) );
  DFFX1 \_right3_reg[30]  ( .D(n145), .CLK(clock), .Q(_right3[30]) );
  DFFX1 \_right3_reg[29]  ( .D(n146), .CLK(clock), .Q(_right3[29]) );
  DFFX1 \_right3_reg[28]  ( .D(n147), .CLK(clock), .Q(_right3[28]) );
  DFFX1 \_right3_reg[27]  ( .D(n148), .CLK(clock), .Q(_right3[27]) );
  DFFX1 \_right3_reg[26]  ( .D(n149), .CLK(clock), .Q(_right3[26]) );
  DFFX1 \_right3_reg[25]  ( .D(n150), .CLK(clock), .Q(_right3[25]) );
  DFFX1 \_right3_reg[24]  ( .D(n151), .CLK(clock), .Q(_right3[24]) );
  DFFX1 \_right3_reg[23]  ( .D(n152), .CLK(clock), .Q(_right3[23]) );
  DFFX1 \_right3_reg[22]  ( .D(n153), .CLK(clock), .Q(_right3[22]) );
  DFFX1 \_right3_reg[21]  ( .D(n154), .CLK(clock), .Q(_right3[21]) );
  DFFX1 \_right3_reg[20]  ( .D(n155), .CLK(clock), .Q(_right3[20]) );
  DFFX1 \_right3_reg[19]  ( .D(n156), .CLK(clock), .Q(_right3[19]) );
  DFFX1 \_right3_reg[18]  ( .D(n157), .CLK(clock), .Q(_right3[18]) );
  DFFX1 \_right3_reg[17]  ( .D(n158), .CLK(clock), .Q(_right3[17]) );
  DFFX1 \_right3_reg[16]  ( .D(n159), .CLK(clock), .Q(_right3[16]) );
  DFFX1 \_right3_reg[15]  ( .D(n160), .CLK(clock), .Q(_right3[15]) );
  DFFX1 \_right3_reg[14]  ( .D(n161), .CLK(clock), .Q(_right3[14]) );
  DFFX1 \_right3_reg[13]  ( .D(n162), .CLK(clock), .Q(_right3[13]) );
  DFFX1 \_right3_reg[12]  ( .D(n163), .CLK(clock), .Q(_right3[12]) );
  DFFX1 \_right3_reg[11]  ( .D(n164), .CLK(clock), .Q(_right3[11]) );
  DFFX1 \_right3_reg[10]  ( .D(n165), .CLK(clock), .Q(_right3[10]) );
  DFFX1 \_right3_reg[9]  ( .D(n166), .CLK(clock), .Q(_right3[9]) );
  DFFX1 \_right3_reg[8]  ( .D(n167), .CLK(clock), .Q(_right3[8]) );
  DFFX1 \_right3_reg[7]  ( .D(n168), .CLK(clock), .Q(_right3[7]) );
  DFFX1 \_right3_reg[6]  ( .D(n169), .CLK(clock), .Q(_right3[6]) );
  DFFX1 \_right3_reg[5]  ( .D(n170), .CLK(clock), .Q(_right3[5]) );
  DFFX1 \betterNeighborCount_buf_reg[0]  ( .D(n272), .CLK(clock), .Q(
        betterNeighborCount[0]) );
  DFFX1 \betterNeighborCount_buf_reg[1]  ( .D(n271), .CLK(clock), .Q(
        betterNeighborCount[1]) );
  DFFX1 \data_out_buf_reg[15]  ( .D(n225), .CLK(clock), .Q(data_out[15]) );
  DFFX1 \data_out_buf_reg[14]  ( .D(n226), .CLK(clock), .Q(data_out[14]) );
  DFFX1 \data_out_buf_reg[13]  ( .D(n227), .CLK(clock), .Q(data_out[13]) );
  DFFX1 \data_out_buf_reg[12]  ( .D(n228), .CLK(clock), .Q(data_out[12]) );
  DFFX1 \data_out_buf_reg[11]  ( .D(n229), .CLK(clock), .Q(data_out[11]) );
  DFFX1 \data_out_buf_reg[10]  ( .D(n230), .CLK(clock), .Q(data_out[10]) );
  DFFX1 \data_out_buf_reg[9]  ( .D(n231), .CLK(clock), .Q(data_out[9]) );
  DFFX1 \data_out_buf_reg[8]  ( .D(n232), .CLK(clock), .Q(data_out[8]) );
  DFFX1 \data_out_buf_reg[7]  ( .D(n233), .CLK(clock), .Q(data_out[7]) );
  DFFX1 \data_out_buf_reg[6]  ( .D(n234), .CLK(clock), .Q(data_out[6]) );
  DFFX1 \data_out_buf_reg[5]  ( .D(n235), .CLK(clock), .Q(data_out[5]) );
  DFFX1 \data_out_buf_reg[4]  ( .D(n236), .CLK(clock), .Q(data_out[4]) );
  DFFX1 \data_out_buf_reg[3]  ( .D(n237), .CLK(clock), .Q(data_out[3]) );
  DFFX1 \data_out_buf_reg[2]  ( .D(n238), .CLK(clock), .Q(data_out[2]) );
  DFFX1 \data_out_buf_reg[1]  ( .D(n239), .CLK(clock), .Q(data_out[1]) );
  DFFX1 \data_out_buf_reg[0]  ( .D(n240), .CLK(clock), .Q(data_out[0]) );
  DFFX1 \explore_constant_reg[15]  ( .D(n290), .CLK(clock), .Q(n421), .QN(n560) );
  DFFX1 \explore_constant_reg[14]  ( .D(n291), .CLK(clock), .Q(n420), .QN(n561) );
  DFFX1 \explore_constant_reg[13]  ( .D(n292), .CLK(clock), .Q(n419), .QN(n562) );
  DFFX1 \explore_constant_reg[12]  ( .D(n293), .CLK(clock), .Q(n418), .QN(n563) );
  DFFX1 \explore_constant_reg[11]  ( .D(n294), .CLK(clock), .Q(n417), .QN(n564) );
  DFFX1 \explore_constant_reg[10]  ( .D(n295), .CLK(clock), .Q(n416), .QN(n565) );
  DFFX1 \explore_constant_reg[9]  ( .D(n296), .CLK(clock), .Q(n415), .QN(n566)
         );
  DFFX1 \explore_constant_reg[8]  ( .D(n297), .CLK(clock), .Q(n414), .QN(n567)
         );
  DFFX1 \explore_constant_reg[7]  ( .D(n298), .CLK(clock), .Q(n413), .QN(n568)
         );
  DFFX1 \explore_constant_reg[6]  ( .D(n299), .CLK(clock), .Q(n412), .QN(n569)
         );
  DFFX1 \explore_constant_reg[5]  ( .D(n300), .CLK(clock), .Q(n411), .QN(n570)
         );
  DFFX1 \explore_constant_reg[4]  ( .D(n301), .CLK(clock), .Q(n410), .QN(n571)
         );
  DFFX1 \explore_constant_reg[3]  ( .D(n302), .CLK(clock), .Q(n409), .QN(n572)
         );
  DFFX1 \explore_constant_reg[2]  ( .D(n303), .CLK(clock), .Q(n408), .QN(n573)
         );
  DFFX1 \explore_constant_reg[1]  ( .D(n304), .CLK(clock), .Q(n407), .QN(n574)
         );
  DFFX1 \explore_constant_reg[0]  ( .D(n305), .CLK(clock), .Q(n405), .QN(n575)
         );
  DFFX1 \address_count_reg[10]  ( .D(n130), .CLK(clock), .Q(address[10]) );
  DFFX1 \address_count_reg[9]  ( .D(n131), .CLK(clock), .Q(address[9]) );
  DFFX1 \address_count_reg[8]  ( .D(n132), .CLK(clock), .Q(address[8]) );
  DFFX1 \address_count_reg[7]  ( .D(n133), .CLK(clock), .Q(address[7]) );
  DFFX1 \address_count_reg[6]  ( .D(n134), .CLK(clock), .Q(address[6]) );
  DFFX1 \address_count_reg[5]  ( .D(n135), .CLK(clock), .Q(address[5]) );
  DFFX1 \address_count_reg[4]  ( .D(n136), .CLK(clock), .Q(address[4]) );
  DFFX1 \address_count_reg[3]  ( .D(n137), .CLK(clock), .Q(address[3]) );
  DFFX1 \address_count_reg[2]  ( .D(n138), .CLK(clock), .Q(address[2]) );
  DFFX1 \address_count_reg[1]  ( .D(n139), .CLK(clock), .Q(address[1]) );
  DFFX1 \nexthop_buf_reg[15]  ( .D(n113), .CLK(clock), .Q(nexthop[15]) );
  DFFX1 \nexthop_buf_reg[14]  ( .D(n114), .CLK(clock), .Q(nexthop[14]) );
  DFFX1 \nexthop_buf_reg[13]  ( .D(n115), .CLK(clock), .Q(nexthop[13]) );
  DFFX1 \nexthop_buf_reg[12]  ( .D(n116), .CLK(clock), .Q(nexthop[12]) );
  DFFX1 \nexthop_buf_reg[11]  ( .D(n117), .CLK(clock), .Q(nexthop[11]) );
  DFFX1 \nexthop_buf_reg[10]  ( .D(n118), .CLK(clock), .Q(nexthop[10]) );
  DFFX1 \nexthop_buf_reg[9]  ( .D(n119), .CLK(clock), .Q(nexthop[9]) );
  DFFX1 \nexthop_buf_reg[8]  ( .D(n120), .CLK(clock), .Q(nexthop[8]) );
  DFFX1 \nexthop_buf_reg[7]  ( .D(n121), .CLK(clock), .Q(nexthop[7]) );
  DFFX1 \nexthop_buf_reg[5]  ( .D(n123), .CLK(clock), .Q(nexthop[5]) );
  DFFX1 \nexthop_buf_reg[4]  ( .D(n124), .CLK(clock), .Q(nexthop[4]) );
  DFFX1 \nexthop_buf_reg[3]  ( .D(n125), .CLK(clock), .Q(nexthop[3]) );
  DFFX1 \nexthop_buf_reg[2]  ( .D(n126), .CLK(clock), .Q(nexthop[2]) );
  DFFX1 \nexthop_buf_reg[1]  ( .D(n127), .CLK(clock), .Q(nexthop[1]) );
  winnerPolicy_DW01_sub_0 sub_131 ( .A(epsilon_buf), .B(epsilon_step), .CI(
        1'b0), .DIFF({N147, N146, N145, N144, N143, N142, N141, N140, N139, 
        N138, N137, N136, N135, N134, N133, N132}) );
  winnerPolicy_DW02_mult_1 mult_171 ( .A({mybest[15:10], N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235}), .B({1'b1, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .TC(1'b0), .PRODUCT({N229, N228, N227, N226, N225, N224, N223, N222, N221, 
        N220, N219, N218, N217, N216, N215, N214, N213, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14}) );
  winnerPolicy_DW02_mult_0 mult_147 ( .A({mybest[15:10], N244, N243, N242, 
        N241, N240, N239, N238, N237, N236, N235}), .B({1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b0}), .TC(1'b0), .PRODUCT({N195, N194, N193, N192, N191, N190, N189, N188, N187, 
        N186, N185, N184, N183, N182, N181, N180, N179, N178, N177, N176, N175, 
        N174, N173, N172, N171, N170, N169, N168, N167, N166, N165, 
        SYNOPSYS_UNCONNECTED__15}) );
  FADDX1 \add_173/U1_16  ( .A(N214), .B(N236), .CI(\add_173/carry[16] ), .CO(
        \add_173/carry[17] ), .S(N246) );
  FADDX1 \add_173/U1_17  ( .A(N215), .B(N237), .CI(\add_173/carry[17] ), .CO(
        \add_173/carry[18] ), .S(N247) );
  FADDX1 \add_173/U1_18  ( .A(N216), .B(N238), .CI(\add_173/carry[18] ), .CO(
        \add_173/carry[19] ), .S(N248) );
  FADDX1 \add_173/U1_19  ( .A(N217), .B(N239), .CI(\add_173/carry[19] ), .CO(
        \add_173/carry[20] ), .S(N249) );
  FADDX1 \add_173/U1_20  ( .A(N218), .B(N240), .CI(\add_173/carry[20] ), .CO(
        \add_173/carry[21] ), .S(N250) );
  FADDX1 \add_173/U1_21  ( .A(N219), .B(N241), .CI(\add_173/carry[21] ), .CO(
        \add_173/carry[22] ), .S(N251) );
  FADDX1 \add_173/U1_22  ( .A(N220), .B(N242), .CI(\add_173/carry[22] ), .CO(
        \add_173/carry[23] ), .S(N252) );
  FADDX1 \add_173/U1_23  ( .A(N221), .B(N243), .CI(\add_173/carry[23] ), .CO(
        \add_173/carry[24] ), .S(N253) );
  FADDX1 \add_173/U1_24  ( .A(N222), .B(N244), .CI(\add_173/carry[24] ), .CO(
        \add_173/carry[25] ), .S(N254) );
  FADDX1 \add_173/U1_25  ( .A(N223), .B(mybest[10]), .CI(\add_173/carry[25] ), 
        .CO(\add_173/carry[26] ), .S(N255) );
  FADDX1 \add_173/U1_26  ( .A(N224), .B(mybest[11]), .CI(\add_173/carry[26] ), 
        .CO(\add_173/carry[27] ), .S(N256) );
  FADDX1 \add_173/U1_27  ( .A(N225), .B(mybest[12]), .CI(\add_173/carry[27] ), 
        .CO(\add_173/carry[28] ), .S(N257) );
  FADDX1 \add_173/U1_28  ( .A(N226), .B(mybest[13]), .CI(\add_173/carry[28] ), 
        .CO(\add_173/carry[29] ), .S(N258) );
  FADDX1 \add_173/U1_29  ( .A(N227), .B(mybest[14]), .CI(\add_173/carry[29] ), 
        .CO(\add_173/carry[30] ), .S(N259) );
  FADDX1 \add_173/U1_30  ( .A(N228), .B(mybest[15]), .CI(\add_173/carry[30] ), 
        .CO(\add_173/carry[31] ), .S(N260) );
  DFFX1 \_right_reg[0]  ( .D(n306), .CLK(clock), .Q(_right[0]), .QN(n553) );
  DFFX1 \_right3_reg[4]  ( .D(n592), .CLK(clock), .Q(_right3[4]), .QN(n559) );
  DFFX1 \_right3_reg[3]  ( .D(n593), .CLK(clock), .Q(_right3[3]), .QN(n558) );
  DFFX1 \_right3_reg[2]  ( .D(n594), .CLK(clock), .Q(_right3[2]), .QN(n557) );
  DFFX1 \_right3_reg[1]  ( .D(n595), .CLK(clock), .Q(_right3[1]), .QN(n556) );
  DFFX1 \_right3_reg[0]  ( .D(n175), .CLK(clock), .Q(_right3[0]), .QN(n554) );
  DFFX1 \epsilon_buf_reg[15]  ( .D(n274), .CLK(clock), .Q(epsilon_buf[15]), 
        .QN(n576) );
  DFFX1 \epsilon_buf_reg[14]  ( .D(n275), .CLK(clock), .Q(epsilon_buf[14]), 
        .QN(n577) );
  DFFX1 \epsilon_buf_reg[13]  ( .D(n276), .CLK(clock), .Q(epsilon_buf[13]), 
        .QN(n578) );
  DFFX1 \epsilon_buf_reg[12]  ( .D(n277), .CLK(clock), .Q(epsilon_buf[12]), 
        .QN(n579) );
  DFFX1 \epsilon_buf_reg[11]  ( .D(n278), .CLK(clock), .Q(epsilon_buf[11]), 
        .QN(n580) );
  DFFX1 \epsilon_buf_reg[10]  ( .D(n279), .CLK(clock), .Q(epsilon_buf[10]), 
        .QN(n581) );
  DFFX1 \epsilon_buf_reg[9]  ( .D(n280), .CLK(clock), .Q(epsilon_buf[9]), .QN(
        n582) );
  DFFX1 \epsilon_buf_reg[8]  ( .D(n281), .CLK(clock), .Q(epsilon_buf[8]), .QN(
        n583) );
  DFFX1 \epsilon_buf_reg[7]  ( .D(n282), .CLK(clock), .Q(epsilon_buf[7]), .QN(
        n584) );
  DFFX1 \epsilon_buf_reg[6]  ( .D(n283), .CLK(clock), .Q(epsilon_buf[6]), .QN(
        n585) );
  DFFX1 \epsilon_buf_reg[5]  ( .D(n284), .CLK(clock), .Q(epsilon_buf[5]), .QN(
        n586) );
  DFFX1 \epsilon_buf_reg[4]  ( .D(n285), .CLK(clock), .Q(epsilon_buf[4]), .QN(
        n587) );
  DFFX1 \epsilon_buf_reg[3]  ( .D(n286), .CLK(clock), .Q(epsilon_buf[3]), .QN(
        n588) );
  DFFX1 \epsilon_buf_reg[2]  ( .D(n287), .CLK(clock), .Q(epsilon_buf[2]), .QN(
        n589) );
  DFFX1 \epsilon_buf_reg[1]  ( .D(n288), .CLK(clock), .Q(epsilon_buf[1]), .QN(
        n590) );
  DFFX1 \epsilon_buf_reg[0]  ( .D(n289), .CLK(clock), .Q(epsilon_buf[0]), .QN(
        n591) );
  DFFX1 \address_count_reg[0]  ( .D(n140), .CLK(clock), .Q(address[0]), .QN(
        n555) );
  DFFX1 \state_reg[3]  ( .D(N479), .CLK(clock), .Q(state[3]), .QN(n549) );
  DFFX1 \state_reg[0]  ( .D(N476), .CLK(clock), .Q(state[0]), .QN(n526) );
  DFFX1 \state_reg[1]  ( .D(N477), .CLK(clock), .Q(state[1]), .QN(n551) );
  DFFX1 done_winnerPolicy_buf_reg ( .D(n141), .CLK(clock), .Q(
        done_winnerPolicy) );
  DFFX1 \state_reg[2]  ( .D(N478), .CLK(clock), .Q(state[2]), .QN(n544) );
  DFFX1 one_reg ( .D(n176), .CLK(clock), .Q(one) );
  DFFX1 two_reg ( .D(n143), .CLK(clock), .Q(two) );
  DFFX1 three_reg ( .D(n142), .CLK(clock), .Q(three) );
  DFFX1 wr_en_buf_reg ( .D(n224), .CLK(clock), .Q(wr_en) );
  DFFX1 en_rng_buf_reg ( .D(n129), .CLK(clock), .Q(en_rng) );
  DFFX1 \_right_reg[6]  ( .D(n202), .CLK(clock), .Q(_right[6]) );
  DFFX1 \_right_reg[5]  ( .D(n203), .CLK(clock), .Q(_right[5]) );
  DFFX1 \_right_reg[4]  ( .D(n204), .CLK(clock), .Q(_right[4]) );
  DFFX1 \_right_reg[3]  ( .D(n205), .CLK(clock), .Q(_right[3]) );
  DFFX1 \_right_reg[2]  ( .D(n206), .CLK(clock), .Q(_right[2]) );
  DFFX1 \_right_reg[1]  ( .D(n207), .CLK(clock), .Q(_right[1]) );
  DFFX1 \_left_reg[31]  ( .D(n208), .CLK(clock), .Q(_left[31]), .QN(n339) );
  DFFX1 \_left_reg[30]  ( .D(n209), .CLK(clock), .Q(_left[30]), .QN(n368) );
  DFFX1 \_left_reg[29]  ( .D(n210), .CLK(clock), .Q(_left[29]), .QN(n369) );
  DFFX1 \_left_reg[28]  ( .D(n211), .CLK(clock), .Q(_left[28]), .QN(n340) );
  DFFX1 \_left_reg[27]  ( .D(n212), .CLK(clock), .Q(_left[27]), .QN(n370) );
  DFFX1 \_left_reg[26]  ( .D(n213), .CLK(clock), .Q(_left[26]), .QN(n341) );
  DFFX1 \_left_reg[25]  ( .D(n214), .CLK(clock), .Q(_left[25]), .QN(n342) );
  DFFX1 \_left_reg[24]  ( .D(n215), .CLK(clock), .Q(_left[24]), .QN(n371) );
  DFFX1 \_left_reg[23]  ( .D(n216), .CLK(clock), .Q(_left[23]), .QN(n372) );
  DFFX1 \_left_reg[22]  ( .D(n217), .CLK(clock), .Q(_left[22]), .QN(n343) );
  DFFX1 \_left_reg[21]  ( .D(n218), .CLK(clock), .Q(_left[21]), .QN(n373) );
  DFFX1 \_left_reg[20]  ( .D(n219), .CLK(clock), .Q(_left[20]), .QN(n374) );
  DFFX1 \_left_reg[19]  ( .D(n220), .CLK(clock), .Q(_left[19]), .QN(n344) );
  DFFX1 \_left_reg[18]  ( .D(n221), .CLK(clock), .Q(_left[18]), .QN(n375) );
  DFFX1 \_left_reg[17]  ( .D(n222), .CLK(clock), .Q(_left[17]), .QN(n376) );
  DFFX1 \_left_reg[16]  ( .D(n223), .CLK(clock), .Q(_left[16]), .QN(n345) );
  DFFX1 \nexthop_buf_reg[6]  ( .D(n122), .CLK(clock), .Q(nexthop[6]) );
  DFFX1 \nexthop_buf_reg[0]  ( .D(n128), .CLK(clock), .Q(nexthop[0]) );
  DFFX1 start_rngAddress_buf_reg ( .D(n241), .CLK(clock), .Q(start_rngAddress)
         );
  DFFX1 \which_buf_reg[15]  ( .D(n242), .CLK(clock), .Q(which[15]) );
  DFFX1 \which_buf_reg[14]  ( .D(n243), .CLK(clock), .Q(which[14]) );
  DFFX1 \which_buf_reg[13]  ( .D(n244), .CLK(clock), .Q(which[13]) );
  DFFX1 \which_buf_reg[12]  ( .D(n245), .CLK(clock), .Q(which[12]) );
  DFFX1 \which_buf_reg[11]  ( .D(n246), .CLK(clock), .Q(which[11]) );
  DFFX1 \which_buf_reg[10]  ( .D(n247), .CLK(clock), .Q(which[10]) );
  DFFX1 \which_buf_reg[9]  ( .D(n248), .CLK(clock), .Q(which[9]) );
  DFFX1 \which_buf_reg[8]  ( .D(n249), .CLK(clock), .Q(which[8]) );
  DFFX1 \which_buf_reg[7]  ( .D(n250), .CLK(clock), .Q(which[7]) );
  DFFX1 \which_buf_reg[6]  ( .D(n251), .CLK(clock), .Q(which[6]) );
  DFFX1 \which_buf_reg[5]  ( .D(n252), .CLK(clock), .Q(which[5]) );
  DFFX1 \which_buf_reg[4]  ( .D(n253), .CLK(clock), .Q(which[4]) );
  DFFX1 \which_buf_reg[3]  ( .D(n254), .CLK(clock), .Q(which[3]) );
  DFFX1 \which_buf_reg[2]  ( .D(n255), .CLK(clock), .Q(which[2]) );
  DFFX1 \which_buf_reg[1]  ( .D(n256), .CLK(clock), .Q(which[1]) );
  DFFX1 \which_buf_reg[0]  ( .D(n273), .CLK(clock), .Q(which[0]) );
  DFFX1 \betterNeighborCount_buf_reg[15]  ( .D(n257), .CLK(clock), .Q(
        betterNeighborCount[15]) );
  DFFX1 \betterNeighborCount_buf_reg[14]  ( .D(n258), .CLK(clock), .Q(
        betterNeighborCount[14]) );
  DFFX1 \betterNeighborCount_buf_reg[13]  ( .D(n259), .CLK(clock), .Q(
        betterNeighborCount[13]) );
  DFFX1 \betterNeighborCount_buf_reg[12]  ( .D(n260), .CLK(clock), .Q(
        betterNeighborCount[12]) );
  DFFX1 \betterNeighborCount_buf_reg[11]  ( .D(n261), .CLK(clock), .Q(
        betterNeighborCount[11]) );
  DFFX1 \betterNeighborCount_buf_reg[10]  ( .D(n262), .CLK(clock), .Q(
        betterNeighborCount[10]) );
  DFFX1 \betterNeighborCount_buf_reg[9]  ( .D(n263), .CLK(clock), .Q(
        betterNeighborCount[9]) );
  DFFX1 \betterNeighborCount_buf_reg[8]  ( .D(n264), .CLK(clock), .Q(
        betterNeighborCount[8]) );
  DFFX1 \betterNeighborCount_buf_reg[7]  ( .D(n265), .CLK(clock), .Q(
        betterNeighborCount[7]) );
  DFFX1 \betterNeighborCount_buf_reg[6]  ( .D(n266), .CLK(clock), .Q(
        betterNeighborCount[6]) );
  DFFX1 \betterNeighborCount_buf_reg[5]  ( .D(n267), .CLK(clock), .Q(
        betterNeighborCount[5]) );
  DFFX1 \betterNeighborCount_buf_reg[4]  ( .D(n268), .CLK(clock), .Q(
        betterNeighborCount[4]) );
  DFFX1 \betterNeighborCount_buf_reg[3]  ( .D(n269), .CLK(clock), .Q(
        betterNeighborCount[3]) );
  DFFX1 \betterNeighborCount_buf_reg[2]  ( .D(n270), .CLK(clock), .Q(
        betterNeighborCount[2]) );
  OR2X1 U316 ( .IN1(n456), .IN2(n427), .Q(n307) );
  OR2X1 U317 ( .IN1(n433), .IN2(n427), .Q(n308) );
  INVX0 U318 ( .INP(n403), .ZN(n313) );
  INVX0 U319 ( .INP(n403), .ZN(n312) );
  INVX0 U320 ( .INP(n403), .ZN(n311) );
  INVX0 U321 ( .INP(n402), .ZN(n461) );
  INVX0 U322 ( .INP(n432), .ZN(n429) );
  INVX0 U323 ( .INP(n472), .ZN(n473) );
  INVX0 U324 ( .INP(n307), .ZN(n314) );
  INVX0 U325 ( .INP(n307), .ZN(n315) );
  INVX0 U326 ( .INP(n307), .ZN(n316) );
  INVX0 U327 ( .INP(n308), .ZN(n309) );
  INVX0 U328 ( .INP(n308), .ZN(n310) );
  NOR2X0 U329 ( .IN1(n483), .IN2(n427), .QN(n406) );
  NOR2X0 U330 ( .IN1(n426), .IN2(n427), .QN(n425) );
  NOR2X0 U331 ( .IN1(n463), .IN2(n427), .QN(n462) );
  NOR2X0 U332 ( .IN1(n490), .IN2(n423), .QN(n434) );
  INVX0 U333 ( .INP(n438), .ZN(n493) );
  NOR2X0 U334 ( .IN1(n422), .IN2(n423), .QN(n404) );
  NOR2X0 U335 ( .IN1(n428), .IN2(n423), .QN(n424) );
  INVX0 U336 ( .INP(n489), .ZN(n495) );
  AOI221X1 U337 ( .IN1(n436), .IN2(n437), .IN3(n576), .IN4(epsilon_step[15]), 
        .IN5(n438), .QN(n435) );
  AND3X1 U338 ( .IN1(n491), .IN2(n489), .IN3(nrst), .Q(n494) );
  INVX0 U339 ( .INP(rng_address[2]), .ZN(N121) );
  INVX0 U340 ( .INP(MY_NODE_ID[1]), .ZN(n400) );
  INVX0 U341 ( .INP(MY_NODE_ID[0]), .ZN(n399) );
  INVX0 U342 ( .INP(nrst), .ZN(n427) );
  INVX0 U343 ( .INP(bestneighborID[1]), .ZN(n401) );
  XNOR2X1 U344 ( .IN1(rng_address[9]), .IN2(\add_121/carry[10] ), .Q(N128) );
  OR2X1 U345 ( .IN1(rng_address[8]), .IN2(\add_121/carry[9] ), .Q(
        \add_121/carry[10] ) );
  XNOR2X1 U346 ( .IN1(\add_121/carry[9] ), .IN2(rng_address[8]), .Q(N127) );
  AND2X1 U347 ( .IN1(\add_121/carry[8] ), .IN2(rng_address[7]), .Q(
        \add_121/carry[9] ) );
  XOR2X1 U348 ( .IN1(rng_address[7]), .IN2(\add_121/carry[8] ), .Q(N126) );
  AND2X1 U349 ( .IN1(\add_121/carry[7] ), .IN2(rng_address[6]), .Q(
        \add_121/carry[8] ) );
  XOR2X1 U350 ( .IN1(rng_address[6]), .IN2(\add_121/carry[7] ), .Q(N125) );
  OR2X1 U351 ( .IN1(rng_address[5]), .IN2(\add_121/carry[6] ), .Q(
        \add_121/carry[7] ) );
  XNOR2X1 U352 ( .IN1(\add_121/carry[6] ), .IN2(rng_address[5]), .Q(N124) );
  OR2X1 U353 ( .IN1(rng_address[4]), .IN2(\add_121/carry[5] ), .Q(
        \add_121/carry[6] ) );
  XNOR2X1 U354 ( .IN1(\add_121/carry[5] ), .IN2(rng_address[4]), .Q(N123) );
  AND2X1 U355 ( .IN1(rng_address[2]), .IN2(rng_address[3]), .Q(
        \add_121/carry[5] ) );
  XOR2X1 U356 ( .IN1(rng_address[3]), .IN2(rng_address[2]), .Q(N122) );
  XOR2X1 U357 ( .IN1(\add_173/carry[31] ), .IN2(N229), .Q(N261) );
  AND2X1 U358 ( .IN1(N213), .IN2(N235), .Q(\add_173/carry[16] ) );
  XOR2X1 U359 ( .IN1(N235), .IN2(N213), .Q(N245) );
  AND2X1 U360 ( .IN1(n345), .IN2(_right[16]), .Q(n317) );
  NOR4X0 U361 ( .IN1(_right[11]), .IN2(_right[10]), .IN3(_right[0]), .IN4(n317), .QN(n322) );
  NOR4X0 U362 ( .IN1(_right[15]), .IN2(_right[14]), .IN3(_right[13]), .IN4(
        _right[12]), .QN(n321) );
  NOR4X0 U363 ( .IN1(_right[4]), .IN2(_right[3]), .IN3(_right[2]), .IN4(
        _right[1]), .QN(n320) );
  OR2X1 U364 ( .IN1(_right[6]), .IN2(_right[5]), .Q(n318) );
  NOR4X0 U365 ( .IN1(n318), .IN2(_right[7]), .IN3(_right[9]), .IN4(_right[8]), 
        .QN(n319) );
  NAND4X0 U366 ( .IN1(n322), .IN2(n321), .IN3(n320), .IN4(n319), .QN(n323) );
  OA221X1 U367 ( .IN1(_right[17]), .IN2(n376), .IN3(_right[16]), .IN4(n345), 
        .IN5(n323), .Q(n324) );
  AO221X1 U368 ( .IN1(_right[17]), .IN2(n376), .IN3(_right[18]), .IN4(n375), 
        .IN5(n324), .Q(n325) );
  OA221X1 U369 ( .IN1(_right[19]), .IN2(n344), .IN3(_right[18]), .IN4(n375), 
        .IN5(n325), .Q(n326) );
  AO221X1 U370 ( .IN1(_right[19]), .IN2(n344), .IN3(_right[20]), .IN4(n374), 
        .IN5(n326), .Q(n327) );
  OA221X1 U371 ( .IN1(_right[21]), .IN2(n373), .IN3(_right[20]), .IN4(n374), 
        .IN5(n327), .Q(n328) );
  AO221X1 U372 ( .IN1(_right[21]), .IN2(n373), .IN3(_right[22]), .IN4(n343), 
        .IN5(n328), .Q(n329) );
  OA221X1 U373 ( .IN1(_right[23]), .IN2(n372), .IN3(_right[22]), .IN4(n343), 
        .IN5(n329), .Q(n330) );
  AO221X1 U374 ( .IN1(_right[23]), .IN2(n372), .IN3(_right[24]), .IN4(n371), 
        .IN5(n330), .Q(n331) );
  OA221X1 U375 ( .IN1(_right[25]), .IN2(n342), .IN3(_right[24]), .IN4(n371), 
        .IN5(n331), .Q(n332) );
  AO221X1 U376 ( .IN1(_right[25]), .IN2(n342), .IN3(_right[26]), .IN4(n341), 
        .IN5(n332), .Q(n333) );
  OA221X1 U377 ( .IN1(_right[27]), .IN2(n370), .IN3(_right[26]), .IN4(n341), 
        .IN5(n333), .Q(n334) );
  AO221X1 U378 ( .IN1(_right[27]), .IN2(n370), .IN3(_right[28]), .IN4(n340), 
        .IN5(n334), .Q(n335) );
  OA221X1 U379 ( .IN1(_right[29]), .IN2(n369), .IN3(_right[28]), .IN4(n340), 
        .IN5(n335), .Q(n336) );
  AO221X1 U380 ( .IN1(_right[29]), .IN2(n369), .IN3(_right[30]), .IN4(n368), 
        .IN5(n336), .Q(n337) );
  OA221X1 U381 ( .IN1(_right[31]), .IN2(n339), .IN3(_right[30]), .IN4(n368), 
        .IN5(n337), .Q(n338) );
  AO21X1 U382 ( .IN1(_right[31]), .IN2(n339), .IN3(n338), .Q(N196) );
  AND2X1 U383 ( .IN1(n345), .IN2(_right3[16]), .Q(n346) );
  NOR4X0 U384 ( .IN1(_right3[11]), .IN2(_right3[10]), .IN3(_right3[0]), .IN4(
        n346), .QN(n351) );
  NOR4X0 U385 ( .IN1(_right3[15]), .IN2(_right3[14]), .IN3(_right3[13]), .IN4(
        _right3[12]), .QN(n350) );
  NOR4X0 U386 ( .IN1(_right3[4]), .IN2(_right3[3]), .IN3(_right3[2]), .IN4(
        _right3[1]), .QN(n349) );
  OR2X1 U387 ( .IN1(_right3[6]), .IN2(_right3[5]), .Q(n347) );
  NOR4X0 U388 ( .IN1(n347), .IN2(_right3[7]), .IN3(_right3[9]), .IN4(
        _right3[8]), .QN(n348) );
  NAND4X0 U389 ( .IN1(n351), .IN2(n350), .IN3(n349), .IN4(n348), .QN(n352) );
  OA221X1 U390 ( .IN1(_right3[17]), .IN2(n376), .IN3(_right3[16]), .IN4(n345), 
        .IN5(n352), .Q(n353) );
  AO221X1 U391 ( .IN1(_right3[17]), .IN2(n376), .IN3(_right3[18]), .IN4(n375), 
        .IN5(n353), .Q(n354) );
  OA221X1 U392 ( .IN1(_right3[19]), .IN2(n344), .IN3(_right3[18]), .IN4(n375), 
        .IN5(n354), .Q(n355) );
  AO221X1 U393 ( .IN1(_right3[19]), .IN2(n344), .IN3(_right3[20]), .IN4(n374), 
        .IN5(n355), .Q(n356) );
  OA221X1 U394 ( .IN1(_right3[21]), .IN2(n373), .IN3(_right3[20]), .IN4(n374), 
        .IN5(n356), .Q(n357) );
  AO221X1 U395 ( .IN1(_right3[21]), .IN2(n373), .IN3(_right3[22]), .IN4(n343), 
        .IN5(n357), .Q(n358) );
  OA221X1 U396 ( .IN1(_right3[23]), .IN2(n372), .IN3(_right3[22]), .IN4(n343), 
        .IN5(n358), .Q(n359) );
  AO221X1 U397 ( .IN1(_right3[23]), .IN2(n372), .IN3(_right3[24]), .IN4(n371), 
        .IN5(n359), .Q(n360) );
  OA221X1 U398 ( .IN1(_right3[25]), .IN2(n342), .IN3(_right3[24]), .IN4(n371), 
        .IN5(n360), .Q(n361) );
  AO221X1 U399 ( .IN1(_right3[25]), .IN2(n342), .IN3(_right3[26]), .IN4(n341), 
        .IN5(n361), .Q(n362) );
  OA221X1 U400 ( .IN1(_right3[27]), .IN2(n370), .IN3(_right3[26]), .IN4(n341), 
        .IN5(n362), .Q(n363) );
  AO221X1 U401 ( .IN1(_right3[27]), .IN2(n370), .IN3(_right3[28]), .IN4(n340), 
        .IN5(n363), .Q(n364) );
  OA221X1 U402 ( .IN1(_right3[29]), .IN2(n369), .IN3(_right3[28]), .IN4(n340), 
        .IN5(n364), .Q(n365) );
  AO221X1 U403 ( .IN1(_right3[29]), .IN2(n369), .IN3(_right3[30]), .IN4(n368), 
        .IN5(n365), .Q(n366) );
  OA221X1 U404 ( .IN1(_right3[31]), .IN2(n339), .IN3(_right3[30]), .IN4(n368), 
        .IN5(n366), .Q(n367) );
  AO21X1 U405 ( .IN1(_right3[31]), .IN2(n339), .IN3(n367), .Q(N262) );
  XOR2X1 U406 ( .IN1(MY_NODE_ID[15]), .IN2(bestneighborID[15]), .Q(n382) );
  XOR2X1 U407 ( .IN1(MY_NODE_ID[2]), .IN2(bestneighborID[2]), .Q(n381) );
  NOR2X0 U408 ( .IN1(n399), .IN2(bestneighborID[0]), .QN(n377) );
  OA22X1 U409 ( .IN1(MY_NODE_ID[1]), .IN2(n377), .IN3(n377), .IN4(n401), .Q(
        n380) );
  AND2X1 U410 ( .IN1(bestneighborID[0]), .IN2(n399), .Q(n378) );
  OA22X1 U411 ( .IN1(n378), .IN2(n400), .IN3(bestneighborID[1]), .IN4(n378), 
        .Q(n379) );
  OR4X1 U412 ( .IN1(n382), .IN2(n381), .IN3(n380), .IN4(n379), .Q(n398) );
  XNOR2X1 U413 ( .IN1(MY_NODE_ID[6]), .IN2(bestneighborID[6]), .Q(n386) );
  XNOR2X1 U414 ( .IN1(MY_NODE_ID[5]), .IN2(bestneighborID[5]), .Q(n385) );
  XNOR2X1 U415 ( .IN1(MY_NODE_ID[4]), .IN2(bestneighborID[4]), .Q(n384) );
  XNOR2X1 U416 ( .IN1(MY_NODE_ID[3]), .IN2(bestneighborID[3]), .Q(n383) );
  NAND4X0 U417 ( .IN1(n386), .IN2(n385), .IN3(n384), .IN4(n383), .QN(n397) );
  XNOR2X1 U418 ( .IN1(MY_NODE_ID[10]), .IN2(bestneighborID[10]), .Q(n390) );
  XNOR2X1 U419 ( .IN1(MY_NODE_ID[9]), .IN2(bestneighborID[9]), .Q(n389) );
  XNOR2X1 U420 ( .IN1(MY_NODE_ID[8]), .IN2(bestneighborID[8]), .Q(n388) );
  XNOR2X1 U421 ( .IN1(MY_NODE_ID[7]), .IN2(bestneighborID[7]), .Q(n387) );
  NAND4X0 U422 ( .IN1(n390), .IN2(n389), .IN3(n388), .IN4(n387), .QN(n396) );
  XNOR2X1 U423 ( .IN1(MY_NODE_ID[14]), .IN2(bestneighborID[14]), .Q(n394) );
  XNOR2X1 U424 ( .IN1(MY_NODE_ID[13]), .IN2(bestneighborID[13]), .Q(n393) );
  XNOR2X1 U425 ( .IN1(MY_NODE_ID[12]), .IN2(bestneighborID[12]), .Q(n392) );
  XNOR2X1 U426 ( .IN1(MY_NODE_ID[11]), .IN2(bestneighborID[11]), .Q(n391) );
  NAND4X0 U427 ( .IN1(n394), .IN2(n393), .IN3(n392), .IN4(n391), .QN(n395) );
  NOR4X0 U428 ( .IN1(n398), .IN2(n397), .IN3(n396), .IN4(n395), .QN(N263) );
  NOR2X0 U429 ( .IN1(n559), .IN2(n402), .QN(n592) );
  NOR2X0 U430 ( .IN1(n558), .IN2(n402), .QN(n593) );
  NOR2X0 U431 ( .IN1(n557), .IN2(n402), .QN(n594) );
  NOR2X0 U432 ( .IN1(n556), .IN2(n402), .QN(n595) );
  NOR2X0 U433 ( .IN1(n553), .IN2(n403), .QN(n306) );
  AO22X1 U434 ( .IN1(n404), .IN2(n405), .IN3(rng_out_4bit[0]), .IN4(n406), .Q(
        n305) );
  AO22X1 U435 ( .IN1(n404), .IN2(n407), .IN3(rng_out_4bit[1]), .IN4(n406), .Q(
        n304) );
  AO22X1 U436 ( .IN1(n404), .IN2(n408), .IN3(rng_out_4bit[2]), .IN4(n406), .Q(
        n303) );
  AO22X1 U437 ( .IN1(n404), .IN2(n409), .IN3(rng_out_4bit[3]), .IN4(n406), .Q(
        n302) );
  AO22X1 U438 ( .IN1(n404), .IN2(n410), .IN3(rng_out_4bit[4]), .IN4(n406), .Q(
        n301) );
  AO22X1 U439 ( .IN1(n404), .IN2(n411), .IN3(rng_out_4bit[5]), .IN4(n406), .Q(
        n300) );
  AO22X1 U440 ( .IN1(n404), .IN2(n412), .IN3(rng_out_4bit[6]), .IN4(n406), .Q(
        n299) );
  AO22X1 U441 ( .IN1(n404), .IN2(n413), .IN3(rng_out_4bit[7]), .IN4(n406), .Q(
        n298) );
  AO22X1 U442 ( .IN1(n404), .IN2(n414), .IN3(rng_out_4bit[8]), .IN4(n406), .Q(
        n297) );
  AO22X1 U443 ( .IN1(n404), .IN2(n415), .IN3(rng_out_4bit[9]), .IN4(n406), .Q(
        n296) );
  AO22X1 U444 ( .IN1(n404), .IN2(n416), .IN3(rng_out_4bit[10]), .IN4(n406), 
        .Q(n295) );
  AO22X1 U445 ( .IN1(n404), .IN2(n417), .IN3(rng_out_4bit[11]), .IN4(n406), 
        .Q(n294) );
  AO22X1 U446 ( .IN1(n404), .IN2(n418), .IN3(rng_out_4bit[12]), .IN4(n406), 
        .Q(n293) );
  AO22X1 U447 ( .IN1(n404), .IN2(n419), .IN3(rng_out_4bit[13]), .IN4(n406), 
        .Q(n292) );
  AO22X1 U448 ( .IN1(n404), .IN2(n420), .IN3(rng_out_4bit[14]), .IN4(n406), 
        .Q(n291) );
  AO22X1 U449 ( .IN1(n404), .IN2(n421), .IN3(rng_out_4bit[15]), .IN4(n406), 
        .Q(n290) );
  AO22X1 U450 ( .IN1(n424), .IN2(epsilon_buf[0]), .IN3(data_in[0]), .IN4(n425), 
        .Q(n289) );
  AO22X1 U451 ( .IN1(n424), .IN2(epsilon_buf[1]), .IN3(data_in[1]), .IN4(n425), 
        .Q(n288) );
  AO22X1 U452 ( .IN1(n424), .IN2(epsilon_buf[2]), .IN3(data_in[2]), .IN4(n425), 
        .Q(n287) );
  AO22X1 U453 ( .IN1(n424), .IN2(epsilon_buf[3]), .IN3(data_in[3]), .IN4(n425), 
        .Q(n286) );
  AO22X1 U454 ( .IN1(n424), .IN2(epsilon_buf[4]), .IN3(data_in[4]), .IN4(n425), 
        .Q(n285) );
  AO22X1 U455 ( .IN1(n424), .IN2(epsilon_buf[5]), .IN3(data_in[5]), .IN4(n425), 
        .Q(n284) );
  AO22X1 U456 ( .IN1(n424), .IN2(epsilon_buf[6]), .IN3(data_in[6]), .IN4(n425), 
        .Q(n283) );
  AO22X1 U457 ( .IN1(n424), .IN2(epsilon_buf[7]), .IN3(data_in[7]), .IN4(n425), 
        .Q(n282) );
  AO22X1 U458 ( .IN1(n424), .IN2(epsilon_buf[8]), .IN3(data_in[8]), .IN4(n425), 
        .Q(n281) );
  AO22X1 U459 ( .IN1(n424), .IN2(epsilon_buf[9]), .IN3(data_in[9]), .IN4(n425), 
        .Q(n280) );
  AO22X1 U460 ( .IN1(n424), .IN2(epsilon_buf[10]), .IN3(data_in[10]), .IN4(
        n425), .Q(n279) );
  AO22X1 U461 ( .IN1(n424), .IN2(epsilon_buf[11]), .IN3(data_in[11]), .IN4(
        n425), .Q(n278) );
  AO22X1 U462 ( .IN1(n424), .IN2(epsilon_buf[12]), .IN3(data_in[12]), .IN4(
        n425), .Q(n277) );
  AO22X1 U463 ( .IN1(n424), .IN2(epsilon_buf[13]), .IN3(data_in[13]), .IN4(
        n425), .Q(n276) );
  AO22X1 U464 ( .IN1(n424), .IN2(epsilon_buf[14]), .IN3(data_in[14]), .IN4(
        n425), .Q(n275) );
  AO22X1 U465 ( .IN1(n424), .IN2(epsilon_buf[15]), .IN3(data_in[15]), .IN4(
        n425), .Q(n274) );
  AO22X1 U466 ( .IN1(which[0]), .IN2(n429), .IN3(n310), .IN4(rng_out_4bit[0]), 
        .Q(n273) );
  AO22X1 U467 ( .IN1(n429), .IN2(betterNeighborCount[0]), .IN3(n309), .IN4(
        data_in[0]), .Q(n272) );
  AO22X1 U468 ( .IN1(n429), .IN2(betterNeighborCount[1]), .IN3(n310), .IN4(
        data_in[1]), .Q(n271) );
  AO22X1 U469 ( .IN1(n429), .IN2(betterNeighborCount[2]), .IN3(n309), .IN4(
        data_in[2]), .Q(n270) );
  AO22X1 U470 ( .IN1(n429), .IN2(betterNeighborCount[3]), .IN3(n310), .IN4(
        data_in[3]), .Q(n269) );
  AO22X1 U471 ( .IN1(n429), .IN2(betterNeighborCount[4]), .IN3(n309), .IN4(
        data_in[4]), .Q(n268) );
  AO22X1 U472 ( .IN1(n429), .IN2(betterNeighborCount[5]), .IN3(n310), .IN4(
        data_in[5]), .Q(n267) );
  AO22X1 U473 ( .IN1(n429), .IN2(betterNeighborCount[6]), .IN3(n309), .IN4(
        data_in[6]), .Q(n266) );
  AO22X1 U474 ( .IN1(n429), .IN2(betterNeighborCount[7]), .IN3(n310), .IN4(
        data_in[7]), .Q(n265) );
  AO22X1 U475 ( .IN1(n429), .IN2(betterNeighborCount[8]), .IN3(n310), .IN4(
        data_in[8]), .Q(n264) );
  AO22X1 U476 ( .IN1(n429), .IN2(betterNeighborCount[9]), .IN3(n310), .IN4(
        data_in[9]), .Q(n263) );
  AO22X1 U477 ( .IN1(n429), .IN2(betterNeighborCount[10]), .IN3(n310), .IN4(
        data_in[10]), .Q(n262) );
  AO22X1 U478 ( .IN1(n429), .IN2(betterNeighborCount[11]), .IN3(n310), .IN4(
        data_in[11]), .Q(n261) );
  AO22X1 U479 ( .IN1(n429), .IN2(betterNeighborCount[12]), .IN3(n310), .IN4(
        data_in[12]), .Q(n260) );
  AO22X1 U480 ( .IN1(n429), .IN2(betterNeighborCount[13]), .IN3(n310), .IN4(
        data_in[13]), .Q(n259) );
  AO22X1 U481 ( .IN1(n429), .IN2(betterNeighborCount[14]), .IN3(n310), .IN4(
        data_in[14]), .Q(n258) );
  AO22X1 U482 ( .IN1(n429), .IN2(betterNeighborCount[15]), .IN3(n310), .IN4(
        data_in[15]), .Q(n257) );
  AO22X1 U483 ( .IN1(which[1]), .IN2(n429), .IN3(n310), .IN4(rng_out_4bit[1]), 
        .Q(n256) );
  AO22X1 U484 ( .IN1(which[2]), .IN2(n429), .IN3(n310), .IN4(rng_out_4bit[2]), 
        .Q(n255) );
  AO22X1 U485 ( .IN1(which[3]), .IN2(n429), .IN3(n310), .IN4(rng_out_4bit[3]), 
        .Q(n254) );
  AO22X1 U486 ( .IN1(which[4]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[4]), 
        .Q(n253) );
  AO22X1 U487 ( .IN1(which[5]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[5]), 
        .Q(n252) );
  AO22X1 U488 ( .IN1(which[6]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[6]), 
        .Q(n251) );
  AO22X1 U489 ( .IN1(which[7]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[7]), 
        .Q(n250) );
  AO22X1 U490 ( .IN1(which[8]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[8]), 
        .Q(n249) );
  AO22X1 U491 ( .IN1(which[9]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[9]), 
        .Q(n248) );
  AO22X1 U492 ( .IN1(which[10]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[10]), .Q(n247) );
  AO22X1 U493 ( .IN1(which[11]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[11]), .Q(n246) );
  AO22X1 U494 ( .IN1(which[12]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[12]), .Q(n245) );
  AO22X1 U495 ( .IN1(which[13]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[13]), .Q(n244) );
  AO22X1 U496 ( .IN1(which[14]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[14]), .Q(n243) );
  AO22X1 U497 ( .IN1(which[15]), .IN2(n429), .IN3(n309), .IN4(rng_out_4bit[15]), .Q(n242) );
  NAND2X0 U498 ( .IN1(n308), .IN2(n430), .QN(n241) );
  NAND3X0 U499 ( .IN1(n429), .IN2(n431), .IN3(start_rngAddress), .QN(n430) );
  AO22X1 U500 ( .IN1(n434), .IN2(data_out[0]), .IN3(N132), .IN4(n435), .Q(n240) );
  AO22X1 U501 ( .IN1(n434), .IN2(data_out[1]), .IN3(N133), .IN4(n435), .Q(n239) );
  AO22X1 U502 ( .IN1(n434), .IN2(data_out[2]), .IN3(N134), .IN4(n435), .Q(n238) );
  AO22X1 U503 ( .IN1(n434), .IN2(data_out[3]), .IN3(N135), .IN4(n435), .Q(n237) );
  AO22X1 U504 ( .IN1(n434), .IN2(data_out[4]), .IN3(N136), .IN4(n435), .Q(n236) );
  AO22X1 U505 ( .IN1(n434), .IN2(data_out[5]), .IN3(N137), .IN4(n435), .Q(n235) );
  AO22X1 U506 ( .IN1(n434), .IN2(data_out[6]), .IN3(N138), .IN4(n435), .Q(n234) );
  AO22X1 U507 ( .IN1(n434), .IN2(data_out[7]), .IN3(N139), .IN4(n435), .Q(n233) );
  AO22X1 U508 ( .IN1(n434), .IN2(data_out[8]), .IN3(N140), .IN4(n435), .Q(n232) );
  AO22X1 U509 ( .IN1(n434), .IN2(data_out[9]), .IN3(N141), .IN4(n435), .Q(n231) );
  AO22X1 U510 ( .IN1(n434), .IN2(data_out[10]), .IN3(N142), .IN4(n435), .Q(
        n230) );
  AO22X1 U511 ( .IN1(n434), .IN2(data_out[11]), .IN3(N143), .IN4(n435), .Q(
        n229) );
  AO22X1 U512 ( .IN1(n434), .IN2(data_out[12]), .IN3(N144), .IN4(n435), .Q(
        n228) );
  AO22X1 U513 ( .IN1(n434), .IN2(data_out[13]), .IN3(N145), .IN4(n435), .Q(
        n227) );
  AO22X1 U514 ( .IN1(n434), .IN2(data_out[14]), .IN3(N146), .IN4(n435), .Q(
        n226) );
  AO22X1 U515 ( .IN1(n434), .IN2(data_out[15]), .IN3(N147), .IN4(n435), .Q(
        n225) );
  OR2X1 U516 ( .IN1(n576), .IN2(epsilon_step[15]), .Q(n437) );
  AO21X1 U517 ( .IN1(n577), .IN2(epsilon_step[14]), .IN3(n439), .Q(n436) );
  OA221X1 U518 ( .IN1(epsilon_step[13]), .IN2(n578), .IN3(epsilon_step[14]), 
        .IN4(n577), .IN5(n440), .Q(n439) );
  AO221X1 U519 ( .IN1(n579), .IN2(epsilon_step[12]), .IN3(n578), .IN4(
        epsilon_step[13]), .IN5(n441), .Q(n440) );
  OA221X1 U520 ( .IN1(epsilon_step[11]), .IN2(n580), .IN3(epsilon_step[12]), 
        .IN4(n579), .IN5(n442), .Q(n441) );
  AO221X1 U521 ( .IN1(n581), .IN2(epsilon_step[10]), .IN3(n580), .IN4(
        epsilon_step[11]), .IN5(n443), .Q(n442) );
  OA221X1 U522 ( .IN1(epsilon_step[9]), .IN2(n582), .IN3(epsilon_step[10]), 
        .IN4(n581), .IN5(n444), .Q(n443) );
  AO221X1 U523 ( .IN1(n583), .IN2(epsilon_step[8]), .IN3(n582), .IN4(
        epsilon_step[9]), .IN5(n445), .Q(n444) );
  OA221X1 U524 ( .IN1(epsilon_step[7]), .IN2(n584), .IN3(epsilon_step[8]), 
        .IN4(n583), .IN5(n446), .Q(n445) );
  AO221X1 U525 ( .IN1(n585), .IN2(epsilon_step[6]), .IN3(n584), .IN4(
        epsilon_step[7]), .IN5(n447), .Q(n446) );
  OA221X1 U526 ( .IN1(epsilon_step[5]), .IN2(n586), .IN3(epsilon_step[6]), 
        .IN4(n585), .IN5(n448), .Q(n447) );
  AO221X1 U527 ( .IN1(n587), .IN2(epsilon_step[4]), .IN3(n586), .IN4(
        epsilon_step[5]), .IN5(n449), .Q(n448) );
  OA221X1 U528 ( .IN1(epsilon_step[3]), .IN2(n588), .IN3(epsilon_step[4]), 
        .IN4(n587), .IN5(n450), .Q(n449) );
  AO222X1 U529 ( .IN1(epsilon_step[2]), .IN2(n451), .IN3(n589), .IN4(n452), 
        .IN5(n588), .IN6(epsilon_step[3]), .Q(n450) );
  OR2X1 U530 ( .IN1(n451), .IN2(epsilon_step[2]), .Q(n452) );
  AO22X1 U531 ( .IN1(n590), .IN2(epsilon_step[1]), .IN3(n453), .IN4(n591), .Q(
        n451) );
  OA21X1 U532 ( .IN1(epsilon_step[1]), .IN2(n590), .IN3(epsilon_step[0]), .Q(
        n453) );
  NAND2X0 U533 ( .IN1(n438), .IN2(n454), .QN(n224) );
  NAND3X0 U534 ( .IN1(n434), .IN2(n455), .IN3(wr_en), .QN(n454) );
  AO22X1 U535 ( .IN1(n311), .IN2(_left[16]), .IN3(bestvalue[0]), .IN4(n314), 
        .Q(n223) );
  AO22X1 U536 ( .IN1(n311), .IN2(_left[17]), .IN3(bestvalue[1]), .IN4(n315), 
        .Q(n222) );
  AO22X1 U537 ( .IN1(n311), .IN2(_left[18]), .IN3(bestvalue[2]), .IN4(n316), 
        .Q(n221) );
  AO22X1 U538 ( .IN1(n311), .IN2(_left[19]), .IN3(bestvalue[3]), .IN4(n314), 
        .Q(n220) );
  AO22X1 U539 ( .IN1(n311), .IN2(_left[20]), .IN3(bestvalue[4]), .IN4(n315), 
        .Q(n219) );
  AO22X1 U540 ( .IN1(n311), .IN2(_left[21]), .IN3(bestvalue[5]), .IN4(n316), 
        .Q(n218) );
  AO22X1 U541 ( .IN1(n311), .IN2(_left[22]), .IN3(bestvalue[6]), .IN4(n314), 
        .Q(n217) );
  AO22X1 U542 ( .IN1(n311), .IN2(_left[23]), .IN3(bestvalue[7]), .IN4(n315), 
        .Q(n216) );
  AO22X1 U543 ( .IN1(n311), .IN2(_left[24]), .IN3(bestvalue[8]), .IN4(n316), 
        .Q(n215) );
  AO22X1 U544 ( .IN1(n311), .IN2(_left[25]), .IN3(bestvalue[9]), .IN4(n314), 
        .Q(n214) );
  AO22X1 U545 ( .IN1(n311), .IN2(_left[26]), .IN3(bestvalue[10]), .IN4(n315), 
        .Q(n213) );
  AO22X1 U546 ( .IN1(n311), .IN2(_left[27]), .IN3(bestvalue[11]), .IN4(n316), 
        .Q(n212) );
  AO22X1 U547 ( .IN1(n312), .IN2(_left[28]), .IN3(bestvalue[12]), .IN4(n316), 
        .Q(n211) );
  AO22X1 U548 ( .IN1(n312), .IN2(_left[29]), .IN3(bestvalue[13]), .IN4(n316), 
        .Q(n210) );
  AO22X1 U549 ( .IN1(n312), .IN2(_left[30]), .IN3(bestvalue[14]), .IN4(n316), 
        .Q(n209) );
  AO22X1 U550 ( .IN1(n312), .IN2(_left[31]), .IN3(bestvalue[15]), .IN4(n316), 
        .Q(n208) );
  AO22X1 U551 ( .IN1(n312), .IN2(_right[1]), .IN3(N165), .IN4(n316), .Q(n207)
         );
  AO22X1 U552 ( .IN1(n312), .IN2(_right[2]), .IN3(N166), .IN4(n316), .Q(n206)
         );
  AO22X1 U553 ( .IN1(n312), .IN2(_right[3]), .IN3(N167), .IN4(n316), .Q(n205)
         );
  AO22X1 U554 ( .IN1(n312), .IN2(_right[4]), .IN3(N168), .IN4(n316), .Q(n204)
         );
  AO22X1 U555 ( .IN1(n312), .IN2(_right[5]), .IN3(N169), .IN4(n316), .Q(n203)
         );
  AO22X1 U556 ( .IN1(n312), .IN2(_right[6]), .IN3(N170), .IN4(n316), .Q(n202)
         );
  AO22X1 U557 ( .IN1(n312), .IN2(_right[7]), .IN3(N171), .IN4(n316), .Q(n201)
         );
  AO22X1 U558 ( .IN1(n312), .IN2(_right[8]), .IN3(N172), .IN4(n315), .Q(n200)
         );
  AO22X1 U559 ( .IN1(n313), .IN2(_right[9]), .IN3(N173), .IN4(n315), .Q(n199)
         );
  AO22X1 U560 ( .IN1(n313), .IN2(_right[10]), .IN3(N174), .IN4(n315), .Q(n198)
         );
  AO22X1 U561 ( .IN1(n313), .IN2(_right[11]), .IN3(N175), .IN4(n315), .Q(n197)
         );
  AO22X1 U562 ( .IN1(n313), .IN2(_right[12]), .IN3(N176), .IN4(n315), .Q(n196)
         );
  AO22X1 U563 ( .IN1(n313), .IN2(_right[13]), .IN3(N177), .IN4(n315), .Q(n195)
         );
  AO22X1 U564 ( .IN1(n313), .IN2(_right[14]), .IN3(N178), .IN4(n315), .Q(n194)
         );
  AO22X1 U565 ( .IN1(n313), .IN2(_right[15]), .IN3(N179), .IN4(n315), .Q(n193)
         );
  AO22X1 U566 ( .IN1(n313), .IN2(_right[16]), .IN3(N180), .IN4(n315), .Q(n192)
         );
  AO22X1 U567 ( .IN1(n313), .IN2(_right[17]), .IN3(N181), .IN4(n315), .Q(n191)
         );
  AO22X1 U568 ( .IN1(n313), .IN2(_right[18]), .IN3(N182), .IN4(n315), .Q(n190)
         );
  AO22X1 U569 ( .IN1(n313), .IN2(_right[19]), .IN3(N183), .IN4(n315), .Q(n189)
         );
  AO22X1 U570 ( .IN1(n313), .IN2(_right[20]), .IN3(N184), .IN4(n314), .Q(n188)
         );
  AO22X1 U571 ( .IN1(n312), .IN2(_right[21]), .IN3(N185), .IN4(n314), .Q(n187)
         );
  AO22X1 U572 ( .IN1(n313), .IN2(_right[22]), .IN3(N186), .IN4(n314), .Q(n186)
         );
  AO22X1 U573 ( .IN1(n311), .IN2(_right[23]), .IN3(N187), .IN4(n314), .Q(n185)
         );
  AO22X1 U574 ( .IN1(n312), .IN2(_right[24]), .IN3(N188), .IN4(n314), .Q(n184)
         );
  AO22X1 U575 ( .IN1(n313), .IN2(_right[25]), .IN3(N189), .IN4(n314), .Q(n183)
         );
  AO22X1 U576 ( .IN1(n311), .IN2(_right[26]), .IN3(N190), .IN4(n314), .Q(n182)
         );
  AO22X1 U577 ( .IN1(n312), .IN2(_right[27]), .IN3(N191), .IN4(n314), .Q(n181)
         );
  AO22X1 U578 ( .IN1(n313), .IN2(_right[28]), .IN3(N192), .IN4(n314), .Q(n180)
         );
  AO22X1 U579 ( .IN1(n311), .IN2(_right[29]), .IN3(N193), .IN4(n314), .Q(n179)
         );
  AO22X1 U580 ( .IN1(n312), .IN2(_right[30]), .IN3(N194), .IN4(n314), .Q(n178)
         );
  AO22X1 U581 ( .IN1(n313), .IN2(_right[31]), .IN3(N195), .IN4(n314), .Q(n177)
         );
  NAND2X0 U582 ( .IN1(n456), .IN2(n457), .QN(n403) );
  MUX21X1 U583 ( .IN1(n458), .IN2(n459), .S(n460), .Q(n176) );
  NOR2X0 U584 ( .IN1(N196), .IN2(n427), .QN(n459) );
  AND2X1 U585 ( .IN1(n457), .IN2(one), .Q(n458) );
  NOR2X0 U586 ( .IN1(n554), .IN2(n402), .QN(n175) );
  AO22X1 U587 ( .IN1(n461), .IN2(_right3[5]), .IN3(N235), .IN4(n462), .Q(n170)
         );
  AO22X1 U588 ( .IN1(n461), .IN2(_right3[6]), .IN3(N236), .IN4(n462), .Q(n169)
         );
  AO22X1 U589 ( .IN1(n461), .IN2(_right3[7]), .IN3(N237), .IN4(n462), .Q(n168)
         );
  AO22X1 U590 ( .IN1(n461), .IN2(_right3[8]), .IN3(N238), .IN4(n462), .Q(n167)
         );
  AO22X1 U591 ( .IN1(n461), .IN2(_right3[9]), .IN3(N239), .IN4(n462), .Q(n166)
         );
  AO22X1 U592 ( .IN1(n461), .IN2(_right3[10]), .IN3(N240), .IN4(n462), .Q(n165) );
  AO22X1 U593 ( .IN1(n461), .IN2(_right3[11]), .IN3(N241), .IN4(n462), .Q(n164) );
  AO22X1 U594 ( .IN1(n461), .IN2(_right3[12]), .IN3(N242), .IN4(n462), .Q(n163) );
  AO22X1 U595 ( .IN1(n461), .IN2(_right3[13]), .IN3(N243), .IN4(n462), .Q(n162) );
  AO22X1 U596 ( .IN1(n461), .IN2(_right3[14]), .IN3(N244), .IN4(n462), .Q(n161) );
  AO22X1 U597 ( .IN1(n461), .IN2(_right3[15]), .IN3(N245), .IN4(n462), .Q(n160) );
  AO22X1 U598 ( .IN1(n461), .IN2(_right3[16]), .IN3(N246), .IN4(n462), .Q(n159) );
  AO22X1 U599 ( .IN1(n461), .IN2(_right3[17]), .IN3(N247), .IN4(n462), .Q(n158) );
  AO22X1 U600 ( .IN1(n461), .IN2(_right3[18]), .IN3(N248), .IN4(n462), .Q(n157) );
  AO22X1 U601 ( .IN1(n461), .IN2(_right3[19]), .IN3(N249), .IN4(n462), .Q(n156) );
  AO22X1 U602 ( .IN1(n461), .IN2(_right3[20]), .IN3(N250), .IN4(n462), .Q(n155) );
  AO22X1 U603 ( .IN1(n461), .IN2(_right3[21]), .IN3(N251), .IN4(n462), .Q(n154) );
  AO22X1 U604 ( .IN1(n461), .IN2(_right3[22]), .IN3(N252), .IN4(n462), .Q(n153) );
  AO22X1 U605 ( .IN1(n461), .IN2(_right3[23]), .IN3(N253), .IN4(n462), .Q(n152) );
  AO22X1 U606 ( .IN1(n461), .IN2(_right3[24]), .IN3(N254), .IN4(n462), .Q(n151) );
  AO22X1 U607 ( .IN1(n461), .IN2(_right3[25]), .IN3(N255), .IN4(n462), .Q(n150) );
  AO22X1 U608 ( .IN1(n461), .IN2(_right3[26]), .IN3(N256), .IN4(n462), .Q(n149) );
  AO22X1 U609 ( .IN1(n461), .IN2(_right3[27]), .IN3(N257), .IN4(n462), .Q(n148) );
  AO22X1 U610 ( .IN1(n461), .IN2(_right3[28]), .IN3(N258), .IN4(n462), .Q(n147) );
  AO22X1 U611 ( .IN1(n461), .IN2(_right3[29]), .IN3(N259), .IN4(n462), .Q(n146) );
  AO22X1 U612 ( .IN1(n461), .IN2(_right3[30]), .IN3(N260), .IN4(n462), .Q(n145) );
  AO22X1 U613 ( .IN1(n461), .IN2(_right3[31]), .IN3(N261), .IN4(n462), .Q(n144) );
  NAND2X0 U614 ( .IN1(n457), .IN2(n463), .QN(n402) );
  MUX21X1 U615 ( .IN1(n464), .IN2(n465), .S(n466), .Q(n143) );
  AND2X1 U616 ( .IN1(N262), .IN2(nrst), .Q(n465) );
  AND2X1 U617 ( .IN1(n457), .IN2(two), .Q(n464) );
  MUX21X1 U618 ( .IN1(n467), .IN2(n468), .S(n466), .Q(n142) );
  INVX0 U619 ( .INP(n469), .ZN(n466) );
  NOR2X0 U620 ( .IN1(N263), .IN2(n427), .QN(n468) );
  AND2X1 U621 ( .IN1(n457), .IN2(three), .Q(n467) );
  AO22X1 U622 ( .IN1(n470), .IN2(nrst), .IN3(n457), .IN4(done_winnerPolicy), 
        .Q(n141) );
  INVX0 U623 ( .INP(n471), .ZN(n470) );
  NOR2X0 U624 ( .IN1(n555), .IN2(n472), .QN(n140) );
  AO22X1 U625 ( .IN1(n473), .IN2(address[1]), .IN3(N119), .IN4(n474), .Q(n139)
         );
  NAND4X0 U626 ( .IN1(n475), .IN2(n476), .IN3(n477), .IN4(n478), .QN(n138) );
  NAND2X0 U627 ( .IN1(N120), .IN2(n474), .QN(n477) );
  NAND2X0 U628 ( .IN1(n473), .IN2(address[2]), .QN(n476) );
  AO221X1 U629 ( .IN1(N121), .IN2(n474), .IN3(n473), .IN4(address[3]), .IN5(
        n479), .Q(n137) );
  AO22X1 U630 ( .IN1(n473), .IN2(address[4]), .IN3(N122), .IN4(n474), .Q(n136)
         );
  AO22X1 U631 ( .IN1(n473), .IN2(address[5]), .IN3(N123), .IN4(n474), .Q(n135)
         );
  AO22X1 U632 ( .IN1(n473), .IN2(address[6]), .IN3(N124), .IN4(n474), .Q(n134)
         );
  AO221X1 U633 ( .IN1(N125), .IN2(n474), .IN3(n473), .IN4(address[7]), .IN5(
        n479), .Q(n133) );
  AO22X1 U634 ( .IN1(n473), .IN2(address[8]), .IN3(N126), .IN4(n474), .Q(n132)
         );
  AO221X1 U635 ( .IN1(N127), .IN2(n474), .IN3(n473), .IN4(address[9]), .IN5(
        n479), .Q(n131) );
  AO221X1 U636 ( .IN1(N128), .IN2(n474), .IN3(n473), .IN4(address[10]), .IN5(
        n479), .Q(n130) );
  INVX0 U637 ( .INP(n478), .ZN(n479) );
  NAND3X0 U638 ( .IN1(nrst), .IN2(n472), .IN3(n480), .QN(n478) );
  AND3X1 U639 ( .IN1(nrst), .IN2(n472), .IN3(n481), .Q(n474) );
  NAND4X0 U640 ( .IN1(n434), .IN2(n482), .IN3(n431), .IN4(n483), .QN(n472) );
  MUX21X1 U641 ( .IN1(n484), .IN2(en_rng), .S(n485), .Q(n129) );
  NOR3X0 U642 ( .IN1(n486), .IN2(n422), .IN3(n432), .QN(n485) );
  NAND2X0 U643 ( .IN1(n433), .IN2(n457), .QN(n432) );
  INVX0 U644 ( .INP(n423), .ZN(n457) );
  OA21X1 U645 ( .IN1(n487), .IN2(n480), .IN3(nrst), .Q(n484) );
  MUX21X1 U646 ( .IN1(nexthop[0]), .IN2(n488), .S(n489), .Q(n128) );
  AO221X1 U647 ( .IN1(n490), .IN2(data_in[0]), .IN3(besthop[0]), .IN4(n491), 
        .IN5(n492), .Q(n488) );
  AO222X1 U648 ( .IN1(n493), .IN2(data_in[1]), .IN3(besthop[1]), .IN4(n494), 
        .IN5(nexthop[1]), .IN6(n495), .Q(n127) );
  AO222X1 U649 ( .IN1(n493), .IN2(data_in[2]), .IN3(besthop[2]), .IN4(n494), 
        .IN5(nexthop[2]), .IN6(n495), .Q(n126) );
  AO222X1 U650 ( .IN1(n493), .IN2(data_in[3]), .IN3(besthop[3]), .IN4(n494), 
        .IN5(nexthop[3]), .IN6(n495), .Q(n125) );
  AO222X1 U651 ( .IN1(n493), .IN2(data_in[4]), .IN3(besthop[4]), .IN4(n494), 
        .IN5(nexthop[4]), .IN6(n495), .Q(n124) );
  AO222X1 U652 ( .IN1(n493), .IN2(data_in[5]), .IN3(besthop[5]), .IN4(n494), 
        .IN5(nexthop[5]), .IN6(n495), .Q(n123) );
  MUX21X1 U653 ( .IN1(nexthop[6]), .IN2(n496), .S(n489), .Q(n122) );
  AO221X1 U654 ( .IN1(n490), .IN2(data_in[6]), .IN3(besthop[6]), .IN4(n491), 
        .IN5(n492), .Q(n496) );
  AO222X1 U655 ( .IN1(n493), .IN2(data_in[7]), .IN3(besthop[7]), .IN4(n494), 
        .IN5(nexthop[7]), .IN6(n495), .Q(n121) );
  AO222X1 U656 ( .IN1(n493), .IN2(data_in[8]), .IN3(besthop[8]), .IN4(n494), 
        .IN5(nexthop[8]), .IN6(n495), .Q(n120) );
  AO222X1 U657 ( .IN1(n493), .IN2(data_in[9]), .IN3(besthop[9]), .IN4(n494), 
        .IN5(nexthop[9]), .IN6(n495), .Q(n119) );
  AO222X1 U658 ( .IN1(n493), .IN2(data_in[10]), .IN3(besthop[10]), .IN4(n494), 
        .IN5(nexthop[10]), .IN6(n495), .Q(n118) );
  AO222X1 U659 ( .IN1(n493), .IN2(data_in[11]), .IN3(besthop[11]), .IN4(n494), 
        .IN5(nexthop[11]), .IN6(n495), .Q(n117) );
  AO222X1 U660 ( .IN1(n493), .IN2(data_in[12]), .IN3(besthop[12]), .IN4(n494), 
        .IN5(nexthop[12]), .IN6(n495), .Q(n116) );
  AO222X1 U661 ( .IN1(n493), .IN2(data_in[13]), .IN3(besthop[13]), .IN4(n494), 
        .IN5(nexthop[13]), .IN6(n495), .Q(n115) );
  AO222X1 U662 ( .IN1(n493), .IN2(data_in[14]), .IN3(besthop[14]), .IN4(n494), 
        .IN5(nexthop[14]), .IN6(n495), .Q(n114) );
  AO222X1 U663 ( .IN1(n493), .IN2(data_in[15]), .IN3(besthop[15]), .IN4(n494), 
        .IN5(nexthop[15]), .IN6(n495), .Q(n113) );
  NAND3X0 U664 ( .IN1(n497), .IN2(n498), .IN3(n434), .QN(n489) );
  OA21X1 U665 ( .IN1(n427), .IN2(en), .IN3(n492), .Q(n423) );
  AO21X1 U666 ( .IN1(n499), .IN2(n500), .IN3(n427), .Q(n492) );
  NAND4X0 U667 ( .IN1(n501), .IN2(three), .IN3(two), .IN4(one), .QN(n498) );
  NAND2X0 U668 ( .IN1(N196), .IN2(n460), .QN(n497) );
  NAND4X0 U669 ( .IN1(n469), .IN2(n455), .IN3(n502), .IN4(n503), .QN(N479) );
  NOR4X0 U670 ( .IN1(n504), .IN2(n501), .IN3(n505), .IN4(n506), .QN(n503) );
  AND2X1 U671 ( .IN1(n460), .IN2(N196), .Q(n505) );
  INVX0 U672 ( .INP(n507), .ZN(n460) );
  INVX0 U673 ( .INP(n508), .ZN(n501) );
  INVX0 U674 ( .INP(n509), .ZN(n504) );
  AND3X1 U675 ( .IN1(n510), .IN2(n463), .IN3(n483), .Q(n502) );
  NAND2X0 U676 ( .IN1(n511), .IN2(n500), .QN(n463) );
  NAND3X0 U677 ( .IN1(n512), .IN2(n307), .IN3(n475), .QN(N478) );
  NOR2X0 U678 ( .IN1(n406), .IN2(n493), .QN(n475) );
  NAND2X0 U679 ( .IN1(n490), .IN2(nrst), .QN(n438) );
  INVX0 U680 ( .INP(n510), .ZN(n490) );
  NAND2X0 U681 ( .IN1(n487), .IN2(n511), .QN(n510) );
  NAND2X0 U682 ( .IN1(nrst), .IN2(n513), .QN(n512) );
  NAND3X0 U683 ( .IN1(n509), .IN2(n431), .IN3(n514), .QN(n513) );
  NAND2X0 U684 ( .IN1(done_rng_address), .IN2(n481), .QN(n431) );
  NAND4X0 U685 ( .IN1(n455), .IN2(n456), .IN3(n515), .IN4(n516), .QN(N477) );
  NOR2X0 U686 ( .IN1(n517), .IN2(n491), .QN(n516) );
  NAND2X0 U687 ( .IN1(n507), .IN2(n508), .QN(n491) );
  NAND2X0 U688 ( .IN1(n518), .IN2(n499), .QN(n508) );
  INVX0 U689 ( .INP(n486), .ZN(n515) );
  NAND2X0 U690 ( .IN1(n509), .IN2(n482), .QN(n486) );
  NAND2X0 U691 ( .IN1(n480), .IN2(n519), .QN(n482) );
  INVX0 U692 ( .INP(n520), .ZN(n480) );
  NAND3X0 U693 ( .IN1(n487), .IN2(n521), .IN3(start_winnerPolicy), .QN(n509)
         );
  NAND2X0 U694 ( .IN1(n518), .IN2(n511), .QN(n456) );
  NAND2X0 U695 ( .IN1(n487), .IN2(n522), .QN(n455) );
  NAND4X0 U696 ( .IN1(n523), .IN2(n514), .IN3(n524), .IN4(n469), .QN(N476) );
  NAND2X0 U697 ( .IN1(n487), .IN2(n499), .QN(n469) );
  NOR2X0 U698 ( .IN1(state[1]), .IN2(state[0]), .QN(n487) );
  NOR2X0 U699 ( .IN1(n422), .IN2(n428), .QN(n524) );
  INVX0 U700 ( .INP(n426), .ZN(n428) );
  NAND2X0 U701 ( .IN1(n522), .IN2(n518), .QN(n426) );
  INVX0 U702 ( .INP(n483), .ZN(n422) );
  NAND2X0 U703 ( .IN1(n525), .IN2(n522), .QN(n483) );
  OA22X1 U704 ( .IN1(n507), .IN2(N196), .IN3(n519), .IN4(n520), .Q(n514) );
  NAND2X0 U705 ( .IN1(n521), .IN2(n518), .QN(n520) );
  NOR2X0 U706 ( .IN1(n526), .IN2(state[1]), .QN(n518) );
  AO21X1 U707 ( .IN1(n560), .IN2(epsilon_buf[15]), .IN3(n527), .Q(n519) );
  OA22X1 U708 ( .IN1(n560), .IN2(epsilon_buf[15]), .IN3(n528), .IN4(n529), .Q(
        n527) );
  NOR2X0 U709 ( .IN1(n577), .IN2(n420), .QN(n529) );
  OA221X1 U710 ( .IN1(n562), .IN2(epsilon_buf[13]), .IN3(n561), .IN4(
        epsilon_buf[14]), .IN5(n530), .Q(n528) );
  AO221X1 U711 ( .IN1(n563), .IN2(epsilon_buf[12]), .IN3(n562), .IN4(
        epsilon_buf[13]), .IN5(n531), .Q(n530) );
  OA221X1 U712 ( .IN1(n564), .IN2(epsilon_buf[11]), .IN3(n563), .IN4(
        epsilon_buf[12]), .IN5(n532), .Q(n531) );
  AO221X1 U713 ( .IN1(n565), .IN2(epsilon_buf[10]), .IN3(n564), .IN4(
        epsilon_buf[11]), .IN5(n533), .Q(n532) );
  OA221X1 U714 ( .IN1(n566), .IN2(epsilon_buf[9]), .IN3(n565), .IN4(
        epsilon_buf[10]), .IN5(n534), .Q(n533) );
  AO221X1 U715 ( .IN1(n567), .IN2(epsilon_buf[8]), .IN3(n566), .IN4(
        epsilon_buf[9]), .IN5(n535), .Q(n534) );
  OA221X1 U716 ( .IN1(n568), .IN2(epsilon_buf[7]), .IN3(n567), .IN4(
        epsilon_buf[8]), .IN5(n536), .Q(n535) );
  AO221X1 U717 ( .IN1(n569), .IN2(epsilon_buf[6]), .IN3(n568), .IN4(
        epsilon_buf[7]), .IN5(n537), .Q(n536) );
  OA221X1 U718 ( .IN1(n570), .IN2(epsilon_buf[5]), .IN3(n569), .IN4(
        epsilon_buf[6]), .IN5(n538), .Q(n537) );
  AO221X1 U719 ( .IN1(n571), .IN2(epsilon_buf[4]), .IN3(n570), .IN4(
        epsilon_buf[5]), .IN5(n539), .Q(n538) );
  OA221X1 U720 ( .IN1(n572), .IN2(epsilon_buf[3]), .IN3(n571), .IN4(
        epsilon_buf[4]), .IN5(n540), .Q(n539) );
  AO222X1 U721 ( .IN1(n541), .IN2(epsilon_buf[2]), .IN3(n573), .IN4(n542), 
        .IN5(n572), .IN6(epsilon_buf[3]), .Q(n540) );
  OR2X1 U722 ( .IN1(n541), .IN2(epsilon_buf[2]), .Q(n542) );
  AO22X1 U723 ( .IN1(n574), .IN2(epsilon_buf[1]), .IN3(n543), .IN4(n575), .Q(
        n541) );
  OA21X1 U724 ( .IN1(n574), .IN2(epsilon_buf[1]), .IN3(epsilon_buf[0]), .Q(
        n543) );
  NAND2X0 U725 ( .IN1(n525), .IN2(n511), .QN(n507) );
  NOR2X0 U726 ( .IN1(n544), .IN2(state[3]), .QN(n511) );
  INVX0 U727 ( .INP(n517), .ZN(n523) );
  NAND3X0 U728 ( .IN1(n545), .IN2(n433), .IN3(n546), .QN(n517) );
  INVX0 U729 ( .INP(n506), .ZN(n546) );
  NAND4X0 U730 ( .IN1(nrst), .IN2(n547), .IN3(n548), .IN4(n471), .QN(n506) );
  NAND2X0 U731 ( .IN1(n525), .IN2(n499), .QN(n471) );
  NAND2X0 U732 ( .IN1(n522), .IN2(n500), .QN(n548) );
  NOR2X0 U733 ( .IN1(n549), .IN2(n544), .QN(n522) );
  NAND3X0 U734 ( .IN1(n500), .IN2(n550), .IN3(n499), .QN(n547) );
  NOR2X0 U735 ( .IN1(n549), .IN2(state[2]), .QN(n499) );
  INVX0 U736 ( .INP(en), .ZN(n550) );
  NAND2X0 U737 ( .IN1(n521), .IN2(n525), .QN(n433) );
  NOR2X0 U738 ( .IN1(n551), .IN2(state[0]), .QN(n525) );
  NAND2X0 U739 ( .IN1(n481), .IN2(n552), .QN(n545) );
  INVX0 U740 ( .INP(done_rng_address), .ZN(n552) );
  AND2X1 U741 ( .IN1(n521), .IN2(n500), .Q(n481) );
  NOR2X0 U742 ( .IN1(n551), .IN2(n526), .QN(n500) );
  NOR2X0 U743 ( .IN1(state[3]), .IN2(state[2]), .QN(n521) );
endmodule

